MPQ    O�    h�  h                                                                                 WI=��
�.�]���Vm��/��H.r�BlQi&�/�-�F>eK��-��~����W�S,��.:j�9�����/���3���V�H��5��:�#m`�Y��[�x����$�x��Z)w17`S��l���;��
�/-�mۡo�kTKg�ơ�O-9{N[�ɴ{d#�$�z �N��M���@�=����P�/]��ab.�YST�{x�"No�H
vS\9����^�Ώ���qj#���V��� o4$�[�/Ez�f�|c�:�6vE	%�pC�3v{�w�A���k��m�[���9��1cTS��M&�S���#:-����gp� I7���-X ��G� �Ԡ�[��b7��Nj}�z3�tN�S�v����8�޺,��9�34}Tπ	{�+�.��B
캿ud�}6؇Աh?
F�!�[�w�0����}U�������q��ܮ�&����Bi��6=�+�=�������]�C�~ϑ��jU�=��Zָ����wr��~�_� ��:����׵��g��!LU��Y�M�o�(���I��˧��$��C���e�وx�yt����R��eX*�¾���B!�6�j)���!7j��U���J�do���x~B�[Vw-o���ԟG���%m�	�����i�+�=�8�P�Q�L9���)�z��/X�򈘳�R#���bBjV�qy,�Agp�����u&<�5ʸ��9 ��}}��r�=r��ЮMZ�]ʬ3{��2�C��tU�(�5$��͓�Llq��i*��1��^JvM�b�I��D��f��&v�����	��]��ݨ�TUi�#�M.J� �BJ5��wS� ������lȾ ��l�N��k���I<��Aj��clw�6�m �M%!I���k�w�%�Y������h�W�X�Q��--D�όu�"09^�TV��+}Oc��l�m)��`���`Cg*V!�"��ك;��x~:e�\���a^��D�OM=w1���ľ�@�L�/�C�K�q��\p�/ Q6L)h�[Rpz';"Q�v�1(���Qbኑ���L�@���#t���8��o���'-	�uG�f6W&i�re��[���"|��Y	0�W(��V�jլk܁u�7�]��+޿�b���Z�?�Y�v�L�ɾѲ�z&0 ��=G�������§t&u���=|ᓵ�jJWyk����x����[�m�U�ȫHM���`��\��{��&٩�����çp3���vR��?�H��R:��
���L�X1ȴ�S�U�E����e�/����&���"�m�}g�x���.(7%�ٕ8�&4���~�؁�ty!�@�
��nE��*��Y�h� }���v���$�f��o[�*����sex&?pZkH��LE���c��T���&���}�P�{��Y��Q�'�suźF}��A�1x|���Շ���iA�U��x2��gH�����L=lP"߭	�2QH|n�u��0p;���s�9�6��\@�q7S��
1���)	-K�y]ٿ���	��6��_�Av�Z�%s�P��t?nc���|�hpٷ$)�
�V{F!N��l�(yK��حS�e�����&+dk�	��w�M�#c�e���ﲪ���6�]�7��Q�B����8(�D���u�Fh�kw������-��H�@0/���#������F���*����o���!�����Ό�܊C�n�{�$W��E��6������n ��&���M�΋�w�?g*X��^f��RUݥxm�&×����]�a�pp��l����ϓ��d�u��?g�p�Ȧrֹb���7�I/���q��DW�\�H؍�s��%��v����?��Ӓȗ����}�;!�a^��9�X5.��HܥD��ڳ��a{��8A���~`��:�l�i�>����+ա�T�4��S�x*ɟU����x�u��Pgj:Z����qU b�s�M��[���� P�3q���[�\ifw~aؽ���$�VV��>BA��h�H��	��y�L����k4w�ʹի�|M�yP��^�B�E�~Y-PCK�(/�}�N��[������g>�c-}AsE�9�M[A�.T����G�Oz���Mo3FQ[-���`f:qO��}��:�%��Ǖ�6�	V\?��#B��[+꡽P�X�ONI�f;j;���}�0� 3�9�Z��·���v�i��%Ge� )�8���Z�8i�h'Wjh��`��*�%�D&Z��s.���w���3��D���X�۹@�mO�.񤷆����n�gK5�����ZTvgM���NV=Ι�Ğ�t�����]���f��w�%\�Q���j�oY���2����m:,x�o�R||m���%��ɋ���^N�Yߓ�}��rQfv�F9(?����ٹ�2l�EX�$X�*�A5/��l�O�����m��|NZ��&��j�7�d�gE�-�X�6T����-k���Z�o*�$F����J*��y:�N#(��*�R�>�D����
���g+P"��J�'�U�z���Y�eWw�����2#D5�0���,�߀��ށy+bGq?n��ԧf�zw"�]Q6��rç|l�˺i$v���0��2��]J ��O�R7h�>�O=��&[X錓nd���k[>��,;s�ЅQh��I{6k��>��E��*�):����<ցa`hq�S}sp�J�_���ɑ�5�$��&e*�Uf+��_�3���k�M%�m�H��4�R�KʛL)��i!�/�C���%6,���F�ҟ���W8E9���̋�<H"��72���t!
P���M���> �.��j�ft^C�Zg�`̸�j-�>��#����~��޷Bx_�bWT��f��YK�w.b/����{��� ]hȏPmc4��u�����d��Kņ����S_�,�}�o���oƌ}������Ng��Ϊ��b��ƨ�/�ޝ�ub�O�\�O��Nݗ|�h���q�er�E�jŽ��_�Dʲ.���!2ܝ&G����[Uh}BhZ3gd��D�±���ƠH�Ue֞�xZ�Zr����'d�ߍ�N�#�Tc����;��/���e�!7�$ي ���.�"u�Ye�6?�˭-!!&@.N�<7��A"�����1�PwvL�.2�5a��N�
b������JX,��6�=F��Q����m�#��L�b��ǞC�M~�Ck�zI��0���
X�j|��s}a}�Y��{S[N�Ν
�N9��׹�,����q����X��l`ooS���=EuZ0��T�:��4v`3�%6�C�Zu{�[ݪ�5�����)0[�k9��1ބ]S^̇&aV�1�5u3�p�+g+�IR�:܂�cX�F�G-/ߥo�N	(a�����z�N����KYOvSיյ{��٘'�/�3��1o/�	�v�+q��}82�Zkp�x�b�/zH?��!'�N���0fmt�"�}�,U��$5��dS��&��-սb��fE+��,�Tl6���؜��9����y�d������R�����Ĉ�_�L]gEA���jg,�w���{�Uy���H�o��I���+��������W�e5�Uxɵ�t����l��:��=�ۮ
�q"j�\�	�7�׌�*b��!d��S�3ϖј-
�<��
GC(�����#��eỊ�!��H��=�-P�R�L����ʓ�Ӗ�m����(���LQBrqt����A��_���x<r�M�֘��t�����}�$�refr��h�]EIB{��~(���(�n�$mH�F;q��'i��_�^�^�(�N\I����zu.�|~7����<��a�3ZԔ�C�Ud���%(J����|55-�SmM���T���� �g��Sk�`�IW".A��,cGO?6A�򞇽!D�S�a�Mw>?YǑ���h�iuWH��셇-(�����"ɳR^
P�Z�+XIc���:;��w�@(_C"9)!	�-�U;���.G��($��P��P�O�^1�c��9��@�Ј/>뇍���+)�.V���$�6g���K�B;P,ҝb��,����u��:���9��|�e�Ř�^���X�N�3�oGv'�@t	�v��2��<�eVl��(}��������w��E���u"�ֈX��������C�uLM��41�'{Ѿ��z�-����GFq�������t��4�ܑ��A֞=J���W�f��FJ�8�_��;�H�5��.M;��`�4Q\5�n˧1�:�ݡ4Z�ÂL����R2�j�C�M�/ו�^�
&�LI�ȏ��O���L���B�/3?��.ľ�!Am,`J�S �i�\%\�h8��[4�>ˣ9%�x�y�ү���#n�s*�*�Y׈W�[Oү�V�/Т$	�ѠJ��eU���es�j�<Z���*�ED��cf�E��w>����?�6{Ӻ�Y��?Q6rsP�2FF\,�1sP{�r
o�q��i\�Z��@�x~$g�H�ŉL=g���^2�n���d�1;�-�sM7�յ�6�Wl��q�Suq�1�K�)�K�XKz�ڴ��	���m�_ky@A�R�Ԡ��P؄�?�(k�j�Ycpѷ(y
^AsF<�����	�]�K�k�����{�@��+�	����#>���ڂ�E[����e��7m��Z/�x��(���׍�uS���f�)����ⷹ��4ͻ�����#Q�Յ/�rz�ֿѡ�ኇً���Ϝ�����}�v�W�wb��]�X� �6N��MD���r��g�Y)��)�mS��O�����ޓ�]x�4pk3�l�þۊK|�h��Ҷ�K�
���7b�-�2%�/w�爴[�_�K\@&��h{�JG�%=ܔ���j?<��e��9}3d�<��t��5�QHד�D�1�Lv�|����ܫ���~��`:(rsi���]j(��p����40�6�S����_�=��u�jz�jAj��C��
�U{ks���\"^l K+�̷i���i���aSփyV� (�U#A�sߣ�_���y0U(;ЈF��w�4��F|�M�^f�I�BoU�~t&�-��hK�b����x5�Ƒ�����c�%A�7e9��F[��.�Zw��Y��x���o�@�Qv
1�'b'`A�
O4I�W-�%�1���6��V1$�#��#��[f�v��8��J_���k;����0���3���!��Rw{�qjϏIdFG GM)��o�/�?8De.'���p�l�%|9�����zI.���݂#F�w?�3�V�\7���+����9�X�+��b��zU\ޢ���4�U��g�gZ��X-J�?�dO,�����]�I��aՇwV-���V�%*���S��oZ���m���j�+|ן�덣���K�"7��4�>����r�z�A׵?k���&��ԥ@lWi*�a�n�e�*5��	��ՀO6���ޗY��Z���E�4��EVN X"�T���L������N����ִJ�r�y5Ԝ~���/�Y�Dw�k�|���v������'�^zHC�t�e����L��m=ߖO0�{,��y��yF�q����¾f���"���Q1 ����p�7jŉ�\��M��y�Y�X�#-�]E+Y��?�R�=ՎYt=R�[3)	�C�h�o}�V4�4�9s{1[Q�KI���k�t?>*��8\)5S��se\�m#a{�
��C9p��X_�Z�d
$5���ׁpO*��fF�Z��3��k!�����	�|�b�K��)��c!r�Cp�H`�6�lA��XW��#9��H�H�kd7m�֕�-?=_�`��^��>;�u�i]A��Cؖ�����"1���L#�z�y��Y�SL���^�x�1�T�Uw�D�/]/�����F�I 8�u#m�.��ph߇G"F�t�8���M�Ӗ����}R������ؼ ��`��i"3�I���=����n�yn��pF�O ���*�i��|����zNC�&�EW�`��ʯ_6�"��BR�<Ñ��3��nS��DU$AhU�:d{����[�ƍb�A���0T<�1�Z�l���'�c��H5s��ST�֙���˿F�+�+(�`�g7-4ኻ���I=luI�ؓ����_�-��@))�<nq����։+S5�A�+�v��k2���a��s�e�q����r ,6���U���� Wbm��,�Sb����^!-M�U�k��
��1�}��5�7߃.9�a�
�YI�W{.L�N�ڦ
�Zy9�����J�T?�q�������spo�V͑��Ep,V�2f�:w5v{�%��zCo�d{�(3�E���%�#f�[h3_9L�1Y'�S9��&K����z�0�{��.�g�a�ImJ����EX���Ghg�
 �[#�AgaX�N��,�p��*�|S�N�+��Ԗ�Ċ��3�.���O	q�+L��������t�s�释b�?��!BiJ�m�l0A�.|�}�������XxW�R�&�9��8|��쮉+0����W���^���Z����������g���.\�&5����_Q��"�+�� ��������Ua��C��ow1u�Li�����p˷
V܅e��x�u�tpQ8�E�'��<���)$ۉ#���Yj_����7 �z��_�3de�h�.�u��l-��e��`VG�*��N���>����$v��l�ۃW�=��P�s�L�
��1�0�ݑ�ʳ���2��B��Jqo����}6Q���<�����9���x�>:X}�ۙ��NrX~��lj]��{eiǳ�����F(���$v.���q�q8i ���T^��Z�u�I�;���a��7����h}���<����u�ޏ�U_��=XJj�4����5���SH�i��<��8 ��E�kk�Irg�A`�Bc"G6V40�9�-!?2Ͽ�%?w�6^Y����Lh��W��*��K
-#��B��"�W�^%k���$+3�Ic=׶ţj��Mԛ��C�g�!7�LS;e�6�B�ʒ�|��_����OÐ
1�T�Ĵ�u@jt,/y
��8+�Ƨ�o ��i�6��G��$&�M;�VG��ӫ�'R��:�\W
��� ���t>���晾3���.\�o��3'���	��L�\�P�wZ�e�T4��L�ؐ��ϴ�qq����� U��R�u�ZN�S���H���mKѐ�B�O���vI�G?Mz\K쩲�ZG�a<�n����t� �7�|7�=�Ҋ���W/���ю�S`���G�#F��>d�M֗o`��7\�/"�b*M�U"|���:�]H��\�R��>"���P$�%Z�Lħ��jÌ��9
{ۍ�?x/����;V
��@Lm�b��.coä"�%�"�8Ê-4G֣��{�"��y ˛�Ψn���*FʄY���A�:�2�J�$�w��%�:���p�K�en��4hZ}�C�E��E��mcAD��&����!pek{��Y���Q�d4s+�:F��c���1nDV��}��,��iwb��K�_x�&Ng���$P�=b�'�c&�2��Pnʗgߙ?;\��s���P���R�����S0f>1�ה)�+jK�W)OT)�OK	4���a _&�fA�ɿ��P�.F?��v�^�e��G�
L�FW�o�FS�EK\6���{�������+�vu	����#�#�$�i�ཛὂ���7(��K����(�:���u��1�aY��Y1��re��6(�6�o!#�����;;��w�r�f��ᥕ���q������y�ùq�WB��2$��-V��$
 a�E�G7�M��W�m��g�zy���}���0�n�5��Pv��z]5Mpf��lQ��E#C��71�����&�\��0�bq�-��/y��C��z�l\�#��C��ǅ��%�+k�� ?o��>SQ�-�r}�����ӯ
K5d&Hҡ�D8�G��,��{T�.H���`~�9U:×�i�K�bH�]���*�4��%�.fΟ�4���yu�Z�j�W���pU���sZߍ�M$��Y� F��'���ri��VaΆp�T�V̟1t�\A�S���v���vy,l���h�!rw�R��M4M�c�龜~B*�$~�M�-FK�������f��a��Uc�i�A�I�9v�,[��A.��H�,w_�e3�M�)o���Q���]`z�Oo�h��?%헭�KA��s�VL���c#�a[�6�����E����T;}H���&�>3�%������_`�lfQ���G�->)��}��=8�'����� C���R+�5�j.E������R�.3W_<���A�ѽU�#�_}�ڿ����U\����6���P�rgdZ>�s����C�*�L�2��],��\��w�T����ޏ��e��ӵ�D�mp��e��|2���HA������/z��9��Hr�W�<�?j��VOS���6lҬ��<j�נ��5U���^ZOp��a��޲����#�� J����EE�|Xv�TIYI�:�Y�,��e������J`~y0�&��Ϡ���t�bD���WR��[�Z����'7�0z�����eM6݃����w�z&0�0�,hh{�4~�ya�q5V��ȃf7��"A�Q,���OQ>���B�Иz.ȇ��径�]@v���R�3�t�`=�c_[�Փ~��
@[QJ����s6��Q���I��kpo>ev4�)f�)04���e�Ly�a�N��I*p��g_t?����5�\��ܛ+*_ tfaO�UD�3�zk\&Zͣ��[ܽ�#K@��)�R�!��CK҅�$�۰<G��U�cW�~93 �́�H�"�7����H� J���53�n>V�D��o��CBuڥDɢ���д�u�#R=�0����Ry.Y�؇���E�Oq�w�FW/}z��C��O� k�>�%m�Ij�k�퇢O"��LASb�|~���!0��}�Z����&�3��kĝل��������8?�_�kJ�O{C�d�I_|	��U����JE�4�ߙ�_��;�����Wt��c�I�M�%�>U��hPGjdzT�Ӎ�ٱ�)���� �c��lͳZ�$��j�'h��ś�9�TYA%Р�Ŀ��;S�6�[,J7�c	�v�
�d�]uĤ�����#`�-W�@$$K<�˦��Me�F������v���2.��a�it��L���>/����,�"}���/#��4�m�%���^bPG�yT�Mt�4k�&\�)Sd� �� փ�}a�(�YĘ�{	]#N d
G�9��B�o�(�tq��o�@�N�Oo�V-�,�aEk�獗U:2��v���%,wKCJD{7k���}f��B�~�j[#�9(+51��S�+&��z�go�+e`�&��g��I�|�x��X��@G��9��_������QVIN�<k��ܷ&=SM@����ϴ���q�3e���O�	�7+'�������p�n�l��j�?;!�!]�M���0�	i�'}&N���l������+F&�ճ�=��~+kj{��cb��݃�T�����).��MB���i�e��{���N_�?�ݎ��9ƌ`�]���6�1U�B��>��o��G����E����˒u���nek_�x�U�t�0�� S��^Z�3���d!l��V�j�Vg�?77{̨��d�^��	^�(�-@�f���{G�_p�	hQ�Y�u�[ �e�۾�=T��PôQLJp�Z�R�Ky,�c����4/�m��B;�;qj�R���8-����<h�ظ����T�ٝ}���(��r î�%];�C{@�I��־Ea(ϒT$�ޓ��q��i�,��kM^������IΨ?�0n���Ɓ �� &�C�Юj�y4JUZ��^t�J%	���P5#wsS#l�2E'�=�� ㇑�_��k&��I���A۷$c�^56�G���\v!: '���w�o�Y���Z�h�ςW����"1�-�eϝ>�"?^@�Lw�+cx :�>����+@���<C���!:5�#6};@��/w'�-������~O~jz1fA�//C@E8�/�I���+�������`�6��S�
z�gI;Ơ��Ge>�"କ�������r?��ل��������)�Io�'Po	�˜��L���e���ݽ��3K�Ҋ�S/½
������uX-��N�8�<.L���ѫ| ��kj�ݐ1���8z��F����G�q�)��# t������߷�i=M{*��>�W�����wB�n��������y�Mq��`�"Z\땕�\-�p�b�*S��8d2�8�SRh�Ɂ9t�����I�@��L?��E����' ��}\�/����T���m"���	������%�w�8�r�4�� ����=�y������]n�g�*��Y��j�TN��/S�e�2$�/c� S��ۻ����0ei��Pr�Z8�W�`�GE:�c�x�M����)�j�a� {I�Yw�Q�s��F���b��1iXM�(����i�8J��Sfx��'g��
ſ��=]��߾�2��an�X�Z~�;7�Rs�����Y��M�D�'��S�z�1�)z[2Kyv��N���B	���GvH_ᘑA�`>Ԗ��P���?���"wYЕ�5��
�v�Frt���IZ'�KAl��$�����ü��0+�,&	�ju�]#��z�_�{@:�Xgn�7���O�nT"(adM��u����\������-1Gz$ͱØ��:#��хe����)��͌�G/D���Sف��v�R�=)��tB�l�uW������Ho�Na� <��~�Mz�A�h��g;����L���w��><÷�M�TA]���pa�ll�|�� ��&[�W��徦#�pb�uy�(5�/ԅ�����ɕ�5\6A������P%s���|cg?�~͒�`R�H��})/��e���}B5��H��]D���ё�+����K��E~��:^�ki��{�72����4&� �	4)��4�s*Vu��Uaщjk�����Uq޴s5Xګ��_Xu� A)��t0��$i�j/aIW�/0�V?C�A����Y��:u7yGȟ�m��@ wTi�|?DM����KQB��O~��A-�2YK�6	�.`j�0��Q�x��c^D�A�{�9�M�[ҷ".�N��>� ����wod�Q�$���^`�I.O��ܭ�r�%�AǦ��gd�Vg��#Әn[�|�!Tw�@�6�w,
;8�4��V�+p3}K�ĭh]�g���ziG�4�)s��%��8���'�녦[��*�U4��L�.,�xܓ�-�3�V����:��oj�~��%���s��XL�0����QX[�Kk�g^����,�KC�5Ɓ���m��]ǒ��WE�w��ʂ&����a�ӐI_PՂm+W�`�|�d;�������H������.��r"��7se?Ņ�����
FlM��=����X5����0O˦�������\�P�۫����!E���X���T�LX���F�Gԭ�ජ��>s�L�J��y+2�4#�[������DmU�2&ȯQ��!Kz���'��8z�(��� e���n*������t0��,�����}�y|�q�0J�x�	frJ"ܻ�Q'@Z��+��_���-��U܇�vA�Y��];�s�`�iRhIu���=Hԭ[��m��"�L�P�Ws�R2Q�\I�MkK�>����ĳ)+5�)���a��U��0�p�l_U���[c5�(	�7�*�yf|ݫЕ3l�(k��>�T�����U�K� �)��0!h��C&�����ҵi�7����{�WiK�9Nd����wH��m7�8�� ��v}���M;>q+��_���dC}22��-���Om�# �K��OЖ	���P��u�J4%w?iU/��<��S�<� �B�y��m4���fd؇��^ڕEn������|+kg�}� ��Q���k�&H�ٟ���?fn��ٴ�Y!%��o��fn�O��EB�/�|�,��0����E�}?�ڈi_�O�_Vs�rE՝��b�$;L�`�U9�FhK�d�M��H<���G�7�~��؞�׿Z�ﱉ���'u��߾t��T�PT��<�{iͿ��_�ݕV|�7�Q�1]�A�u?zē�m��^��-�7�@?�<$F
�r8�a-ā73���E�v�
�2ɍa�OQ���@�ݙ#	,,���vK�jY��V2m����]�b#ꞔ�%Mkr�=�d�-��Y�kh{m����a�f�Y?��{�.N[S�
��v9�&8�ʯƏ��q�1�'�)��o ����xEf0�����:��v��%��C%�{rͿ�{'3��m��>[�"�9C*#1O��S��&�H+���&ᯁ]�g\gRI�����X�}�G�7��@��� ܿ����s�N�r�fU��MS��=�L�o���@�@oV3 `	��	ga�+:��.���+e�i��@��?�T5!x�Y�c�b0�����&}����@���?���&F��.��"+���%�L��|���7j6F�D������֤���\X��f?_��c��T�ӌ��j�*�qJfUJD��9'o-���G�7D�����m��Fke�Mx�U�t&0^�=	�Ѡ���I�?V�"'ej�.�	
7���A+0�9?�d[/l��=��G�-�@��l}GT����h�t���;��@b���=�.@P�L��t���f|���b-�jjS����B��Dqe��Tv��C{�&n]<�;�g�ާ%Q�t!}�����`rΡF���]��6{a��/�b�O8(�T$,��w? qڑit���o^6�8	PI�56狚���E����s�@��$J�s��vUUu����J�K���5�T�S����mm���ƒ ު���)�k�iWI�Q�AV��cؖ�6�z��o��!5�Z�r`Bwo��Y�[�
Πh���W�͵�6�-h9���"���^[��5t+钄c�IQ��+����N�Q�CS%{!U{i�?�;ߴj�%��[���݆�a>�O9d�1��Ī�\@ �/�L�nrk��?�S6�������4;��I��@��W�	1�	����)�f���ʢ)��$�QoX�'�"	*~�RL����:�e'D�ݸ"��%N�E��۽��!��T�WI�u�ƈI'_��3;�N����D��E7��ˉ��K�z�昩���GW�|��FK�>�-t���m�K��Y�=�CⵔeW���w>��0ٕ�J��G�봜M��`}ɸ\F��حѩ��������'�s��R=��4�^XP�ƽ��["�L�v�� q�� �9�	��x�/Dt߂������m��;��f>��E%-�r8�z�4��K�j���X�,y�v(Cn1@}*|iYȡ��l�쯰����'$zޠ�:���B�- ed7`���Z��ϖ{��E���c�I����=�U�s����UV{Y-�RQ}!�s���F��/�1d�`σ������i�.��A�x�رg4���ZG�=X���H2=/6n :�Ղ?;��s�%ՆP?�Hj����S��1
P�)��fKT���hAڅ�e	>����p_�X�A�E��Pi�W?Z89�;��T0b���!
��3F������5��K|�d���q��؁�Q�+P	��uO�#��!��,4���N��Ѕ7�Czc<��ϝ(<�N� u$���W���Ҿ��n"�(�,�)�_{�#A�� ���Ɣ(�����+�����Q26�x�ъ�W��gV	W�ν���c�l�ɽ� ����=MI��c�Gg���J����%%�d�Ò^����]I��p\��l	ۻ2ݹ�5��I���&1�^+bP���#��//=��<�ɰ�\�~K��w����%+@�w�?%a������c��}��v�����%�5���H��D��5�}@ڑ����$�e�o_�~LV�:�B�i�In���zY��4��'��!�Ag}���u��m�4�j&�9��kU�G�s�֫�l��V <��4�Gg�i��Oa�ω�
t=VB�����A�'�ߴɈ��Y�ybD���ވ�/�w�3��Q�M�͐�Z0$B�D~��^-<}#K[��i5��S����a��ӻ�c?�A�͉9l��[��3.@���b&���ܷorQ�a�䘣,`�9�O�|��(Ž%�ð��B"uuV�<��g#�3�[�����;R~�Ҽ?;�_�	2��3X��F�"�#�r�b���Z6kGQ[)4q���8�ן'C��A��1ݟ�����q.G��������3�m��-Ӌ��Aۤٝ:�as�Hi�ӣ����S	���"�F`g�����|�
���h��&����]bgf�R�mwg��=y�X�[OV�k��!m�j��[�|����ܲ�5 �������> �i �r�P��2q�? C��� "�%��lȓ)��/S�7�5���O&����|<��:Íˠ��e��PztE'p}X�} T�_ðhءb*o�[Ў���⎇�J��y&���ak����;�D���t��d�����2�'�:!zy�����eCũI��L��{;0��,qv���)y���q++�S<�f��|"w�Q" ���9�h
��7esژ0��
���]6l���R#+����=�d�[Ĩ^��n�@%�G��E�vs�4Q�4@I)�k&�>ۢ��_!_)&V(ǄƼ���a̴�?W�p[b5_��ƽ54'5�HגR�*խ#f���K�3G��k�~_��������s�K�b�)e!�a�CJp�N�P2+ �=�W$8�9i�Q�w�cH���7�~i��Ưq���>��{�����;�C���z�ٸ�
崪�}#�"f'��m`����N8��Ie��E'w���/�xC6,�� � �:��Km��H�a��X
��P^1�KT�r���d��e�}#�i�z�w��%a���jٺRѺ����'%Ɣ*��J�{�a��O1�� J��5�|�������Q�E(��՗ _G>��*�6c�������U��MhF��d0g��V���V��^i������ZSa�����'��$�yD��o�TOv��Vc��֗�a�Q��7>"���r�ƚ�8u�o<��T˙�-��@z�<୫-�N�|ʷ��s룼��v8V2d@}a�U
�v�޷���,�i,�t��q����Oamէ�=N�b�S���MjyVkMR�����NU��,�)��_ma��eY��X{���N���
}�I9�i�%�$���q�P:xY��o[%X�b|�Eab��CZv:��v�C�%"�0C 6�{�Ot��w��K�4ۥ[�JF9^I�1���S�S&���❸�!����$Bg�I�^�n)�XgzpG�d��~���ҿRޢ���N�A���F�U�S�f������P�ě�-3�(����	�Dk+݌M�i1ԺƁQ�d�f����?��!�jm����0Ҥ��G�}\�k��4$�ir$�ȇ&�wթ�\�}Iw+�Қ���n��;�
��%���_P����!���iɒ�������_b��SXD�oI�V�?E�3��$�U�e��4|�o����}�x�R���y.}�H��,|e�X{x�u�t�O!�vH0��ù)�]����]9j0&S���71A������T�d� �=ς�g-vz��"[G�*9��3֏ܛ�Qw���4
�=���P���L ��й!����Y�p�E�����Bq1fq`h �Ǯz�A|O<^�B܌�`m�D}���~�r�c����Q]1�u{���j�{^�(�66$�2��2�_q��i��l�x��^q1���SI�����N�hf�6v��E��&�F	�ݯ�;UP���C�J����!�s5R�S�@���c�sT ���� k�WI���A�(Mc��k6ξ�
��!0�j��-Tw*AY3�a�h`�PW4jL�X\c-A	�S�"��^v|	.+�@zc���t���SyԬ��C��!p�>iU;�7|�?��cW���L����O�}�18���%��@��/*(�	ُ�Sŧ�{�����6��� ���;<�_�}�˰�KG��9c�$T�h4Am��J���
/�l�o��,'�k�	E���͡����(�8e���ݳ���� &�8	�� 9"۱���u�2ƈD�a��X��	����,���"T�&R��lz-d㩣�4G��\���5�Y�ct}���H�B�-�=�,���2W@��2%���Q��t������h�M�2x`x�S\�¼˓:���� �9���얮�aR����/x��)�ׁ�Źv��L5����w�;�?L3��s�/�p҂l���^�m*O����U��%Ȁ�8��K4X��%��s`�y��%�Q�Xnl8>*i�YÔn���ʯkK`��d�$� %��B��Q�)���e_�M-Z������!E0�Dc��k���%��]�[��{��pYH�Q���s�Z�F2���Db1_���ޗ�]�i�D�����xy��goM���y=S���t��2���n;�P�1;�<�s942�!g��CT����Sa;1%<%)pK/d ��� &'	�����_W8�A���Ԍ�&PD��?�}�����O�ʷ�e�
J,�F��8�w�8q�K��I�Z/��#����w+�S	
�\�+#�I�Շ�����d�$��7Yľ:��dk(���f�u��$�R���j�	�(=`5ͧp��:1#=����n��a����<y��*�wش�,��γъJ[�b��WS%|c);�~�D:/ ���l�M���^0g񞪺����i;�߭��m����]�agpW�(lb�4�vj���dG�\nӷ������b��%���/�)�t���˙�\,܇�Ԅz�6(�%��>�r�T?�c_�o� �~�3}F����\�`�-55�_HË4DI'��8G��볉��k�J�]~��:��Di��������� \4�:��/��|0Z���)u����Rj��~�+cNUg��s멃��@3� 7��8�����i�a?���זV}�FE�A��4��V��^ey}������>2w�_ղ��M�2��4�B[Բ~��-��yK6�@��*���*������.�nc�Y1A�?�9��[�au.{����-���˷^r�o��Q⾹���`�I�O ����7[%މ��\qݥ�V��!�#���[RR�W��6���-m�;��=�8�33�W��+¾ٟ�]���G��)O����^8��%'~ȅܢR�X���f�.b ��n��n�3����4��3��4ϥ��D�+<f�Nh�0�ގV`��Kb�AŐg3F����\�++������3]�[w�M5�w����C/����\��F�$�e�mA�ـV�|C���y��P�A�ٶ㠦���UrX��-��?{ �����@f�lC7���B*�Q�W5&�խ���O��@���(��1�F�O��#���iE�"X�19TZ�V�k�}�X��	��c���J1�y!.�y���Ŝ�Dc>���-����WÅ�|`'H��z4V���?�e�D�$�8�Y�K]z0��,y%��e�]y�5�q�ED�.�Ff�t�"5�Q��`�g�#Փ�R%���a���E���K�]1���R��%�œ�=>�[�h�/����G�BLU���sg��Q�,bI~$�k`�>i�����)!�@��&�}\�a������p6x�_ˇh��,5� ���݀*��qf�Y�Ƙ-3"]jk[��thu����Ρ�Kq�)4!^>CܵLz�����-ͱ�fuW�DS9��5��%�Hi87Y��Tg�0�����J]�>�)��Ug-��cC��WY��BY��x#�Eu����E+��?�@���t��@�w�/I&�)�̤2	5 �R��\mjY|�\�A��������������?�ქ}��ϐu,��D��������N�5�;�%��S����N�\O��������[�|z�w���j�7�E������_�L����G9��EG�ڢ���W(Uo��hA�!d��SӾ���2�ͩ-޿˜O5�L�Z��4��Y�'+5M�44.��fnT�@�1}�2,�$^�L|�7��B���mƵ�"u5�`�}���� �-(�@՟<ښ��������s�-���svs��2��a�{��ќ���f�GS�,"�Ѩ����%����mИ��^b�:@�ʭ>M�o�k(���v��V��1e{��aC�Y5�[{�OUN�K�
�T9��׀\C�@F�q���؀߷�o�������E\�����:ch�v痭%��EC���{��ݱ�4��9�쏗C[T��9y��1E��S�Ś&7���8����7g��SI�2K�閆XB�PGT�H�v>��f����M�N��\���_S�)}����������d3�����	]H�+��I���^�a6�_އ�C)?l�!�U��Y�0�¢!�}��m��Hf����>Ǟ&9�n�$".�X|+�8�[Fɠ�ǜe���)��zh�|��ӕ��Y��������4_��Qm����&��� �,���U����/�(o����8(��mRj�����#sXB1�e<Ax��6t܎�1s{��s����h��'Aj�=]����7����vc�o�KdQ0���]�Ͻ.-�z���G
�-�:ʺ֪4���V��׺�o0P=%��P�7�L[Q໋�ϙ��I�ԏ�� 6L��B��q[�uc��i�5�\�i<��s��꧛�/���}���9�rrDE����]�7{�ر��L'��(�8�$�sϓ���q9ic>�Sp�^���U�I����AS�#<�Qe8i��HT�f��J�UK���o�YJV1j�<�5�o|S����P��� �PS�p��kWe+I޻!AL��c�f6BAA�`!+*W�(�w���YN¸� �h;�_Wo�?���-:�Ϯ'�"p&�^����+� c)<<�m=����9�C�b�!�g<��;Ѱ���>��r�����O��b1SY3Ġ�s@�C�/e�I��_ۭҧ������6�q��{���s�;w?���ư&w��SC���?]T��^���ӱ�_g��\5o�j'�F�	`�8�H&y#�c��e]��ݮx�D: һ��S&e�{��ی�WͿ�u)e��?@�M�9��pR��4*�;.��n���3سz�&��C�Gc��Z��t��t�L��#��h��=5���2W�/���+6���m1�����*U<MB�@`sw*\��p�N�f���ơ�����w���y�R9�l�**��<�ٹ�j�L��0�֞@�v�9�|�ns�/��ł'5L�4��m���MÐ�E%c5r8��4�cB���s���yy��,�n�P3*���Y��
�"K�&	M���g$p8��j2���d�"�eZӥa��Zi?얱OkE�N�c�ύ������?�
r�A{z�_Yc��Qs^�s���Fm�K3��1ZT��9�χL�i�z��7��xT
�g�]|Ő��=N�����2��+n6\���o;��st�ռ���>^��8IISyW1@H�)�K
�;�)ڻ�`	��^�Xs�_8*A����P�?��ѝq�JPϷF3
�hFúv��3�E K�\c���H���2��{+��	%r|kE#��`�O�L�&ᩚ���7egU�ͬ�&Y(�%u���uZ8f�M�g�����^THXJ�"wo��#xC#�6^��-���Cx��R��)�����~�]d�W���k��z���� ��E�3�MKF�YitgL@{��R���͹�Z���H�t��L][`pR�@l��R�1��	���zӒ
F��e�b�C`��M/���/���Ӏ\�Ypد�r�q�%D���mL�?ۅ�*J�Ι��}�j���5ӛ�!5�6�H�jD�t��������]�%E�~��:/n�i�<8$�ɿIb4�;W:4�GZ��]�����D��u���r[�j��g�FIYU�zgsƂ�95+)� 2�Q�{��z�i~ia��Ӄ�[�V�ܠ���A�{�j��k��y����8��m�w(��M�DM���Y�B��~�)2-2r\Kdt��?;������:bc���A��9bn[c��.����U�}w����o��zQ�;P��,`�y�O[�0�^��%�o$Ƿ,���V�����#d�7[�Ok���N�1�̈=+;i�w*� �L3}d�'��YB��X�r�OG�k)j�E����8�\'�Sąwv���!�f,��!.})���a���J�3C��c06��EѤ� �K;��FP��ɲo����ɸ��"��<�=go�{�(�赔�H��@��B]�p �H�hw2�ʳ~�Jx��Q���!����m�I��Q�m|�{�4���k����Qc�{.G��r�:�(�_?���B2��[&!l���uq׌3�5�P���OܿK�MĘ�q���������ƌ�E]��X��T��E�&�硘6j�Qc�>yю���J��y��E>Hό`���PD��(��a<�������'�m�z�*����Qe94l��f|���C�^10�D2,��q� =�y͌�q!��	0�f#:x"��vQ�/ﻎ��޿��mgS^���A8���%�*#`],��q��R�Jd����=��a[zH(�j�k�v�[=��L�s"�cQ
ElI�?/k��>QO���\�)�T�:�}8�la���5�p�C_y��kE�5�L�H��*K�cf�G�AJ 3�=�kHW5��Y��vl�)x�K,�&)O��!�:�C�A����҆��(����;W�q�9�P��mm�HD>�7������ͯ''��>���������C.*���q���i�`�#>���;������r��h�����;=_wP��/�D 5��1� �k*��m��W���ET������h������;}Y�-�p希����W�H���ѰA��#��
�O��a:�W�kO�hv����|����*��ǋ7E^����C_�z������xW��+���(��sU
Edh<��d����y?��Mڬ��}��w�K�X��Z��*�{>d'��u��Cg��m�TE+���H�m�D�zb�G,�7�`�b�,�з�u��0�X����C-�n1@P4<5u���$I��d���T�r�bv�L�2��a���,���qAA�b�,���_Ǆ���'��m˩��b<v���`�M`��k�B�����������/a�Y�^�{u�pN�a
��9ۻ����!����q'C%�������o�s�͘��EW&y���:E�v�%��C��"{#���L�i��v{��s�[��9��1�3S�W5&rP��ӁV���g��
I�|��d$�X�`G�``���9��#��nN'Q7��~q`S9��`vȻl�Q'�3Qf�	�kO+������]����ZuQ�Q�	?'�}!�`��Ԃ.0� �U�}����|ė�����Y&Tȍ՟�+�3�0+W�����[�����r�Ә��<����)C�Uh}�-�!��d9_��ɡ���l�Ld���"9�U	��*��o>��������	ܭoCB��\}V�e�ўx�Nt7�����"'̹e��дq��W}jfu��*�7�5��rLcъ�Fd�`��u�o��TH-��ܥ��Geu���*��Ŭb�GN�����۪v#=��P��_L�1V�Fq��E��OV��� �YTB��qV`��L�$H	�w��<T ��=���ElP}�N���r�Fj�
J�]'��{��t��G�۷(�Z�$=Պ����qT�i�
|�.w^��,���I����ߟ�,�ltU�
ِ��������UF=��ʑ*J�Q�Wy�5��S��V��p�� �Ӷ��p�k�{I��wA��ci��6}��@�	!&x��(�w���Yi�C�{�h�W�����"-
S��	`�"+j�^���0�+z�cd�Ū=����"�b�yC�1�!�b�;�I�Yʙ�������r��Oj�1n��Aq@���/����?��'<�P�:�L�i6	����mb�;�	ߝ��9�kL�������Z���^�������â��/�loi��'<A	{X�ì/Th�{�e���ݩS�t9�v=ncֽ�ه�g���uķN�:����I��N�]�ɶY��I<3�n�ozc�`���]Gh����Ꮸ�tsñ��T�ߣ��=�]���n W�ꧪ�Rz��ʻ��.�j���ea[M�9A`n~=\Wo��	cW��o͡ŵä�$��R�ب�%��o,R��ҹ�>�L++ȱ具��'�楍i�/Uɸ�����O�}mO�u������%�	�8�Rl4��5�����y~�i��n�\*M��Y��b�}�G���}��n�$�Q�l������R��eU����Z$����ϜE&�c���9mR�&���&ͮ�{5��Y~c�Q�,�srv�F�M8�%91U�Bϔ�)��ʗi��
���9x/Spg��_�+��=IIQ�*�2n�LnQ��FP�;��s����W�`�9�T䓲�S�X1[t�)fY�K�1�vw��V�	��H���_�WeA3��Ԃ��P�_k?h���Ep����
�a9F޼\�ma��:�K-��>H��%�bn�+�C�	@_d�*#`i��K�ڲ�%��ڰ�7�%tp�r�Z�(�p�9��u����H�Ώ 3 ���s�f͝�$���A#�����6����9z
3�>�,���m��� �)Z슀�n�X,W	29�̙�M�:�� �N�n��M��[�T�g�,�{?��R��՜��#��@��]u�pM!�lnp��9c�!#T����m��C�b!�2��p/@#�����.�\"�؊��Ǭ��%ߙd�h/2?6�����δ��}��^�^�֊i5k�H��{D��볮*M�,|��	<� �6~���:�3�iص�j��Vrb4ƅ�u�5��"���,^u�"^��jW��aO�U]D�s�{�tI��#: -�S�m��x4�i#oba5�ꃛ��V���{��A�U>�ŵ��&�#y�x
���h�w@R���E5M�\�k��B�S&~��-��K�]��u��$�F��Q���ucJ�A0��9�c�[>��.��n�3�ExL޷�1oPÜQٮ�	_`c�6O�����|%�u(�ܰSg�V�t�Y#?�[ȥ���
��,e=��-�;$��E��Ů3�"������B�S2��k(1G���)�+��v8fjB'��t�j�����r���ӻ.�r-�d����Fd3~s'������wV��ؓ�a���Dj��^��;뚽�I�7�fg�1��Ą���!Mq7��Y.�]3�a�C��wx�^�n1e�p���e��|�<v4mw�<�L!�|�m���5�Ɇ������V�Ҷ�r�O�#+?1;e���F�v�l9�u��(���&5\ƌ���_O7ע��9<'�<��g���FE���X���TZ���e��죙��[�"Q�8nJJgX�yn_����G�����DY�����X�=rT�el��p3'�6z�W�82e�C^��e���z���`0��E,/��ۼ�y��q��n����f^"H.�Q Z��#���Ӊ����u�����w����]'�z��NRT����=4��[UH����h���8��V�s��Q%}^It{hk���>�U��0*)yeǕG��a�M����p�#_A�h�~5���ףT�*��f�U/��3�>lk�s.ͪ�v��܄n�K�Gy)j�+!TW�C���¨��!�G#q)�A�WU�C9�45��԰H��7�A��O'��j���sr��>ݧJ�K��c�CigZ�K !������#������;�uy �����q�6��w�2�/���_�e�(z� Z�Ye6{m��k�R��iځhڛ�����ǲW F}�փ�k�ӌ��B��}�%��+ 9�_���E���=�R>�OB��1�#�|p������ uE����Ƅ�_X���K����ɽ��\���g�L6�U��sh7)�dAsz�4䭱h��#=��R�R��@yZ$v��vC�'�]�ߪs�����T�5�����6�Z�i�B��7O0��C����u+��3���JA+-^@�<�o�^j,��aC�#��ME�v���25�a�'^��Ǭ�,��}�,|Q�:"x�Vra��hm�ڀN�b�Ѧ� 4xMۼck�e�P�?����;
���6a:��Y+��{P�<NGģ
Np9ւf�6����	qB�x}���O�oK��3XBER���Tn8:�Av�z%���C��{^�J�������Ep[ʁR9�f,1;��S[	�&�=��nu����:$gH��I���ѯX�0�G�X�����,�cu~�*"NB�^�RwL�St���(ȶ*Ĭ��3CM,P	S��+nE���к����U����tj?�c�!�ٴO�0c^��3�}-Q����>�z���$�&o����U��+�ߐ��}&��8˜q)V�<��Y�r���ݤ֐��Ȭ���N�_s�m��a��r���=�o��]s�U����%;&o�Kg®�%���խ��v��f���'er��x��t�m+�(~�=�̹�j�۫i����j͙��u�7B�P�-B�ѥ3	dG��P���3��-Gb��G�J7������D����ϣ��V���j=[%@P��L2L�}����0��<��ց����
BB�ZqQ�B~��ހ��f<�A��Ӟ�����o*}�Ų�!�r�h��%��]��{���;<LJ=(���$�V&�c2�qo*&i�%�	�Y^"�f��.I���������d􁇣�_$�^���a݀KUA��%iJ̖]�r�5�
�SjJ�YN��D�� �v��&s�k��I��ABcD��6��B�ۡ�!!�ÿ�U�w[kOY������[h�}�W�D��)�u-�a�d�"��x^ǭ�zo�+U
�c��w�E.�����Խ�C? �!�ӯ���;��V\(�4
+��Yq��7&O%�'1���Ė�@��/�e�������������6$���q׿HqD;���N%�	Н�\�N���uK�����:m���颕����o��F'�[Z	���>b�/͈�{�e�� ݤNO�β�1�����q���B�C��u_*׈5�����:���2��1��$�K���z�����E�Gã���u��5t�Y��ٺ����=T�����AWQ���c�b��謕y/�E˚렍.Mx�y`i��\�u��4��x�������_ȬRo�<� ���]hײp���2�L���ȌL����	pЍd�/�%�����j��m�ҋP���%���8���4iR��V�ȁ�^gy�����[�n�*�'�Y�-w�؏毜���#�$f� G�l���NeP�[�SZ�0���o�E�uicc�!�tۖ�����?(�-{��Y��Qi�sM4=F�Ƹi��1P�����#��i�iG_�-3x
��g F��Ƶi=D��߅|�2)2nl�k���;~us�R��j�4�~��;PS��<1v�^)�(qK������j<	�Ѯ��_���AN4���ƬP��<?F���a�@����
{,.F������+�O.Kh�2�+�����Ӽ�xC+<��	[laQ�#;)���Y������fw5��7���������(��[tY�u�3��C�1�{����3��������,#���l/{��%���r����G���,���u��d6�&�S�Wd�7�No���҄�o ��&���M����O�g㼺6L.�*��PĲ�����{�n]���pH��lsz�ۧ�B�<�&�xS7�Hn��J@�b�l��0/�Z��a���\��E�ek����E%z���c2;?�*���U��\�}����9����53H��iDZo��ic�9|<�]�۪K~8�:eOi�N�Ԋ����q��4�d��Pa�-Li�z}u��(1jP&�|u�U�-�s|����}7_ߠ (ԑI|Ë3i>��a��M�vÃV.;���A�O�� � ��,Yy�t��܈C+Vw{� ՃםM�!���qB�Cf~1�%-(��K�w�U���������?9�cj�AKV�9Xy�[PZ.,\y���s��oA�o�Q3���e]`>9O�i��OD%ϛ�m���"V�y�Á#�C[��(H��'Vu�>>;��`���3��-2
�s��N�c�G=6Z)�����D8A��'/Lم�}���V�١��.�����Z
�tb�3�
��A���7�E#(���|���A�w%��?��X���2�g%�w�G ��2�L������]��:�>��w����)���ȵGE��י�w.�m���GԬ|T�>몓�ɡ���� �1���UmWr);<���?�xG���pّl���^;P��<5�[\��4"O�p�Ë�T'���X�B��<�E���X��Tk�Ü������Gv���ꀎsRsJ��yMR��%�T���Dԋ��y)E�xa�(<E��''Y �ze4ݶ1�ze/s����Ի
u��0��,�n��\y�qUV����f�$�"��?Q@ �q�T�)��K��� ������`2�]"��'��R���{W=��+[0h2��ǹ��ol3n��W�s�V$Q@�8I�֍k�`�>�{���J)r��?�_Za8 �+1�p�y�_|�ƽ��'5~]��?w*�H4f��7*3�_�k����ES����
�߄ZK�)�)�	!ϓ:Cm���Ҽs�w�gW+�9�8Q�c\MH��7
�֕��2�7ů���{�v>��J��~�>\C����i���^�"+#�mt�ϋ��#@PF��:\��c��1�w�/z�z�^��� 5Z����m;�'�M
S���-�<��K�^�H�������}�Ґf��U�8�ͺ6�&��Ѧ��:��ƀ�P���Y�MsO��\�D6�&�x|�[_�w�A�=�fE��½�V_�7��7���:l���ػk�v�ՆU@2�h2�d���宅��r���L�-\I���IZ�g~�qh0'<"��e�����T;`�����A�	�=�e7�������u��Փ�˅G-�ݠ@��<뉽��S��~W�����(2v$�I2�Jya�������#���,��s��ۗ�H4�]Gm�+b�O!b�M �'!MV+k�)���6����SB���K��aU}�Y��n{+b�N���
���9�i�בO�q�Cq]�0�i�pˠoGB���6EMjr�_9:�^:v8T}%�Cl3{���݂W<��P�젌[�)�9��1�^S6ۚ&�J��	�+5��H�Zg%�I*q�Z�FXӭGq,�G=D�?���G~�N]N�͏�'5RS�3ӵSU�ȱ��BK3ǋ�G�3	��+I��U*��2���P�,�=K?�7�!���ʿ�0>�L�l�}ȱ�|D՗���o��&�DՕ����,�+�#K�,I)��w'�v���������d����恒c���XW_��?k���~0�Bc����ͻUQ,�� �o��:�i�g���W�e�7˴��� �e�"x�5Qt�o�b�5�X�u��iۆ>�I�j�D̙��97�����W/�� �d�!��+}�n+y-�D(��:kG@L�kL����Ʌ=��L� c&=�rlP���LlR»����k��EC���Wz��V�B�S�qL�Kt�Pǚ������<J����&�L�{�<}�\	J��ru�V�@#]�k{b�j�V���(��J$������q��i}�;��,^]:�&�I��L�RXq�T�ց��'�O��9n\2>���@U<���`,J�y����35��SE4m��N�ߔ� �9�����k�N�I/�{A��/c��6�Z��v��!tD�9�\wd+Y���q�h� .W #ӵ�2�- �!Ͽ0�"�Q�^��͎+08�cڗs��>`��#=���C�.�!ܹ%O;b�z�P��υ��H��(UO�$01�l��
Q@goi/e|�u���{#�����u6?F&���#��;(�.��n��Uk���t8U����T�~���6�#�0=���o�'���	����7G
R%��e.��ݟiEUIl��|��=����g~�u��7�0e�^.���s�M]ɬ9���Ծ�Dz������vGt���Q��.�ti��@��`�=��{FW��� ��'ƕ�p� ����ٵM��`d�\��&�����>b�Z�#��nR
6)� 5%�^�m�n��F�L!,d�g��'I��s�_�/���X�h���}m��+ ^�A\%4f8���4����;)��H�yt�]��8�nXYK*���Y��G�3bůW����$�":�"�u�=�툂veK-�r� Z���0�E9�c>���iO�\K��T���{��DY��iQ�)�s(6F`��p1Kpf�J%��I(�i4�����,x�D�g[�B�a�)=?g����&2�_�n�><y�;YL�s%1�Ս0�/<�I�SM�1�,B)\�K��~��-ڌl�	���i�;_C��Ai�`�xGP�S?��͝B�;���W��
6GF!!�cL*|��K�m���o���>��+��	v���!Z#	��4�����;x7E���t�P�(�fw�?Iu+���>`���7⏗����͓J��H�#)���HZ��Qx��y�ה�bx��c�"��V�Ο2؊��չN�oW���O��ꥠ�0l� ^���ɖM���JOjg]�-��x��E����B��0����]PpCrlΦ��b�&�Wa������#P^��]�bW1��
e�/����`J��7B�\�2�@�{�"	�%�j�^U ?쬄�[S�����}(қՠ�L��5��)H��3D���$��T�䉋м����~sM�: �i��5�+�z�ۡ��4#�+��h�����uz
��fj;����jUS7�sW����K��? ##�����biY�,a+6��Q�Vi���
�A�i��{HO���ry�B �i���w�t��~M���!�DBGS�~L��-��LK��p��?��Z�b��������c�AfH�9ӮL[�4\.gܷ�i��n"���o��QNs����'`�O�y�/BB%�������ɨV	����#��[>�o�å��"g�̙n�;�J`{I��Җ3���m��*<F�I��!��G���)�GA�H?8l'j��H����3K�w_+�RWl.�d��Z��O�*3����4�J��;u���|qs�Lk�:9Rp�z�F���-�,g��U2tI0��u�';a�Ϩm]in��9�tw.����r��ȵ���Ӳ���Fm����B�f|��2�enɼ���z1��ڶ�P rą�G?�Չ�s��٬&Vl/��9���=��5�$�}��O��m�~�o2=�2�ȫ[c�w	E.ӥX�A5TƠ��W�M�鸏��/����`��VPJ�ORyL�Vy4Ͻ���1a7DO���T���p�2v���v'�)�z iG�L�+e�����E�;�#'0���,�6�QXyR�q��ɓ���f�I�"~��Q	����L`�@����w�8�w�E�1����i?]g���R�k��1�=*C[�/�_�G�.d��sS�Q[M�IjR�kmK>�A�f%q)�z�K�_iK�aSd����p��_���<Od5y�(�YK�*|�f�a��3��.k�=��6X��4�:��K]+k)�BZ!J��CH��8W^�Wa �����W˷�9�\���VHբ7E���z�${�8lY6�[>���AqE$C�A祁)I��bC�q٦#og����1af+3��u��P���,f6wa׌/5b�o�k� �&�<�mփ��HXf�������٦��-��<�}*��a���������s�A{}�!=g���ƻ8��Qs��H� O�Z����A4	|f��R���xHE/���9_����9��b�yW��F�U�NU�ؚh-��d��!Ӫ�?��S�K0�	�ZZy܉l�P'��� 3+��BT��HН$U�����@�8��7/���A�!N[u!���*w���-���@�Z<Fġ��U���3���v_�'2k�a�S��=r���*��3�,����7���>{���lm��?�bm��6:�Mщ�k�oY�ƻ�U�r������0ap{�Y!C"{S�N��C
�w�9�p���5>�,M?qx��nvˀKg1o�YC�i58EH<y�
q:O�=vS(�%�;�CGX�{ԺH���������Ȼ[@�9���11�TS�e&#x�⤟z�����g�wIE��Ռ�X�J�G@���|�r��zQ9�UNx��HȠ}CS�v���Ȭ��b�3��Gb0�	I�+$���x�ͭy�Kp��b%�?X+k!BJ�E�g0zP�D}c2g�w؇�0���*d&�j���-��up+����4d��ֿ��ͱ̐���Ul�hl1?���V�9���p_)�
���������Y��r��G�U��[�oOT�$����a��҄ˏڨ.��e��Hx��<tH���^�s�ƹ����a3����jj7ܶ��kw7��������d=����ϩƏ-}G�ǐ�GvU��&���م����bC��[	V=���P���Lǒ��w���/8��ix��M��
�Bx,vqG� ����Ul\�Ȣc<�����D����׆}{��.�r0s�[��]�i'{=H�������P(��6$N�����q�ai�������^����nI�#,�D:�4���a�U�^�*mQݶ4�U7%���w]JB|ᆨ'5�%�S �����
�z�� �J��ׄkC�IJ*A8s�c���6.N��7!"���Ow�|kY��T��"�h���W[!��_�-�]���#"\�q^�çpL�+��c��{o���g��s�xC�]n!����v;=Բ�d��j!&��Wϗ��CO���1�]Č3@B�/Q�5��o�U��a�E�}�6Z"�gvT��l;c(E���c�����]K/�������H��;�q�q����\Noz��'m�N	�ʦ�4-U���O�e�[ݚ����eҧb���ڽg;��S�,�u�op�+kS����s��h���'�@���;q\z4�ᩊ��Gyd@�FM����t������T�i=��+�v��W�n�ن�+��o3ݳ�L�F�M���`_S�\h���:8©-뒡��*�5���ՖR��m�2� 5�(���z�L���Bz��b˪S㍍Z��/f>��о���m��r.�|7%�G�8�J�4������R�y�ڛ�5�n��*G&Y�3���T�@��"�J$\�}��I,�x���#�veF��͟MZU�֖�E��c[v��|���x��e�'{f,DY�dSQ_X�s�FYv�g01Fd"ϥ���FiO���#hx��_g��B��,"=:&��;�`2��Hn� Y�=b;4�3s` ��(���*��䤮�S��1���)�'Kv��'�l�'��	�[�Ąd_�v/A����[mP��?�����Z6�����
�!�F/������W��K�]ҭaŗ�~ze�s�+��n	���W�#����/v��R3ᕲ��b7 (���Ѭ�T�(^�EJuƮ�9��1��JC.����ь끞�#d�����Q�ڝV�J|!d6�}���ޯ��sW���N\�QMݹI lW�u
�f������_ 9�G��$M��L�E1g����4�`�ĥFs=ô�u���`]��p>�zl)���a�r0d�n�$��Q1���0b�;�݂/Q)h����R�\�����4�]Q�%�(�Y��?GO.�A���l}�p��,�Ӈ$:5<a�H���D���4E�o|u�d_����~��L:�D�i�����L�5����4�Q�Uh���W��~�uu�K�(;j�Mu��!U�`�s2&5�%F�� ������!pit�a����,��V�RLq�A������}30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��} ��UWP�Hh1�;�f��l݇�Jߚl�.�u?W�������Jd�WT�VEk_+�o�y�wϢ�w�Yc$�����^�l]b���
_��Dd�3ٱ���k	�9%]���^Al����}���V<�
=��s�'KK9�#�~v����B�I<���[�z��!������c��D�P �=�����:����e��$^�]�]��.�(� ݿ�E�o�hO��z�Sp[�(�혾��K�Ǿ)J;ǜ�zH��z: >ߌd����+|�"�<�H��l�
�M�tc��X,�D��e�b)��n+yL(�f7X2E�3�.�/���1��7��؈MsQ������{�+'|�.��C��@�7_����i�)j��{�!� ۷͖ٳ���U�!�0��\���� rbExy��⵭��T�cUc� �'�a6&~lx/~"\�&���+.G�����k/�~��<�Q�]���/�UZ4Dn��&]�\ֲ	0���+e<�6�p����ꓭh����@��#c	��N�
N�p��Z�(��xmW�wyM��({Cn$�]x�I���b
�^_�Izmh� 5X��.��,���$J�K6��\����ᡊ�J,+%��� ��^�����Brn����WwJaÍ���>\�D����Kq�Ţ���c���"��Y�P(�=�q�#�2n��M�I��6
���d��!N_W�q\[���#AC �+�n�K�PDL�������㳙���/t�]X5Q�����K;�?Ч�4���\X�%>��f�$X�9�}���u�I�����I�e��%1���X���ь �v�����]����iC����F�c���{ֿ-�����N�f!Q�\������8�qe�ϱ	}���DT}u�Rf`a~�O�R�a���tI��.>*[�y��t��Tq#f�K��Wxy	����Fa��)����86P�Y}X���ݍ�s�g���zB����R��C��70,�ԍ�h�R��_��I^��g�Ѻ��fH��N��,z �%6�t!u�K�!g�A�l�١�9���/�A�G\s��t��~u;�Kp壓��[.�/�V�Aפ��Io[C���$�z�k4f��8X��W��5��(t���۹�nl\�4W�m$d�,���X�c6Z��(��MeT��+�u��;'�;�:���!�(��+t�(|�d�pFV̢-���ʹ��JS~L �� ���#J�#��A�C,�,�*���S�ӟ��]�� ����mkVQ���^��N<G+#'���b`}������K�V�=o;�WOhVp ��O���f�Q��y�qk�(�6��)2���K�}�뇾�č�C�qռ��B��
����
�Z���}�K`BbOBlN��bWw���D5S
�T�oQ�'�X�p��dÈ��KW|7�\
�֩�+m�Lv�1%fm�"d���	5�u�1O���	x��jOg%E1dIv�Ҷ�VW�^
�j|��f��h�������SP�3/��;/�r�[-�G5�]���k���X&e<a#@�=��4���	��rD�7S�?�x	N����	o���$D��ߞ@�3�r4!�Ť���c�#ӳ��rT[�?ο����`��Ր�P�Q�¡WZ�6T��q���^Ck�=�+&��v��LY��_���rkw$��ʇ
sc�1t��n&\~x䦀8��[WN�F�T��!��ps����Un�p����AM8�g�A�r�����t�y�q�����f��IM� ���RAKkˇJ'j�q����ߚ�?�S������)4�1U�Z'?#�,'��yh(��T���²M�4${a٭<����v���ˎs��ǯ��!F�x=�f��R�x�̳D�J�㎿J�s�������؄�+F��h��q`�p�-��|짽����v��R�1Ŀr��z���dyB;�q#����c1'zݺ��<��_�`���L��B�a6�f��T�� �����!<*�7z�H;�]	�kS� N�OiMe*�k-��^A��.����b��^��W �iD)<�Ԯ�;Ư���|�C�A�DQ�����������H'�:fPs�񿆃C������w�6T�/�P"^��tPa6u�G��_A;+��޸ދ�1��ۯ⧨������c81�k.x�+���_DP���[��s!��%$�x������.I��ň.���:-�w1�����$��)up��^��J�觭��W�I���O"�4�������k�^�[�C�3�p���=xw�*�<Yd�٫L>0!* ���˼h�����	�EL� ^ �{J�Z��s�	�������J��nW��V��&_������Xw��~$�üHl��!��Ha_�ϵd"h�2�~��9���>ulڅH+�Q��K�n�2ƅ/\'!}�9_�e~I�P���?W�a���Ɖ�3��N���Mx��� R���x�����łe>��$q�L�к�.�q; #�E�q�[Kt8�szu�[�&�|"��Zj�~�{���kǏ��Hk��z��ߟ"����+O��o@M�L�����̠i��{X?j�e��b�2ԡ	Syߚ�f*Eݖ?.����$�>��]�s�9��x>�{�3�|m.��9V�n@tf_b	j��[�)�5�{�l� .am�I�ߌ�*KUV����d��+���U��y^?�h���gn�Uy�)�^X'�Y*&k�/q�.�y����G���L~�Q}<���]���/�i4� ���9��oI%	�����@<�������Aح�QV�l������	:��N~��ۣ
Z����k���Qږ@P{V�H���#����f���O�<WohܛR5�=l���i�KKy����~�8`�H��<(����J��0+8W�Vc�1��������O��C��J�����\�����b�~���5+=�	������~(�qP�\2AR����I��f6�� 
l����_j�7qυ_���HC3["���Ku|,Lh��C�|��$���/G8�Xhg��U� K.SB�������\*F#%�1bf�İX���}����'?I�����x�t%�=�+����x�	����M����fɝ��G}�c��h�u^-R�5��	ԜKQ�]�� ��mZ�����g���Z���}}ȅ�fe��bdG��g_s�D�2Ԣ*�.s��2����f��K��bx�~��z��O�Ja*��� ?8�o����<�����:������h �R�3�q���8u�(�$�an�R���_��^��1g�X;�D̮�˳a�%,�ڠ��2tM�I��x�g�Gl� ��K����A��F��t�0�X��>O�D/�"�AJ󭆕�d�J;z�ʗ���ΚQ�����IGZ��(���n:a�c��H�m�+,+O��Z6-E(�M��`��@X	���ZMcI
���M�py���ʹ��^��V]&Pe���~r�i�����3�� �\��ڜ��S������!G��`��S��l�j�h�������n1M�7�6zP�����/��'+K{��v�[Ã1��Dǩ6�&�a�H��gfv+�nip1#􅃢�o�@f������]��4���ؐ��!�1�P"�0'�������ٍd],�!"�"R/{�\.G�f7h3�Q���gO�OC��rs��WDܻ eG�@7M�~<�zI�: ?��۔f��
��D~���IO���^$��&�U*���ы��1V*�Z��_wbS.�����:[���9؃��װT���Po���ÙG�;�Sq�p��=�9���E�Ŧ)	b�6���9>�e�]a��ta(RM�
3��i�9�Њu3痂ȓ�;����z�  5�RLx��,zd}��P��ˈ��#��Z~��B�J0® yC��:����U|Qd�>4�"g>�q�g�yJ�C����K��:��TS4�T�ޒ�)��W[7��W`M��qSu$��"ԥ�:dtj-<�n�#�`K��U+�f3\Q�tX�P0=�J��-����K������yC�ӈ�����L#�����k���+��5p}�����Q�Yq�f�ͱᐓ���b��+��B�1���7�ޢn\�����u�?_&�?��B�2oU��xټw�n��ZS�奀�(�uw��d�[i�uջ��@�&�e)�l*��A���VÚ�J���Z�F'�Q��"�+]���y;Z:�g��(�G���h���Wޏ=��l�vP�	�3ir.�eS�2(��Z�B���-����ؿ"�@]��rE���E,�F*{#}GV�\]���e����
�,���P�G�,2Z�ԁ���q�=�^� *=�
�&�;�	��S����a�ka�b���0s�&t^]&F���+8+�nW�g��>�a!�s.G9���Z�Z�q��%M�����}�\�Y��H�@�q�	E��d��`QM ٨-Z�+��_<'Ԅ��;|w��z�?1��kx�OZ+4|�lU�v'��,�|yR=0���:c;�\'�4����(��.j��m��]8����I6�Fl\��PR��v�6�*��2����s�z<�����rG����h����`~#!-�������JC���	����1�zy����&B%��#���ͥ(z��5��s�����9f��5B�����T0������a����^�U9� x8\i�m�*��)A<�h. �E�=t�H�WJi���~�c;�ģ�/�C9�D��}�|.`�[^V��'}dbP]����0CA�t�l���a��T�pi��m^f�,PK��u���"�A�#A���;�������Q���ք����xH.��pn���T��[D����%Nӗ�+�����lIɒňX��Ѥ�{�!�m^~��B���Yu�	^���{у�X�~�"�"�Y���q��^��AC�&lp'������#Y�@��r�W0�TI��:��z�%�Ƹ���� �D}1J<L'�+����1�@�t�x�5J�w�Wq�VR�_����v&�ll�w�V�$|[g�f��lz����^_�hd�jv���	��9�1�+�kl��U>"�R/0���o��'K"9��~���ݠ�j2�UXP�s�M��} �@b���~ <}�����-Ҙ�,e(��$���:�t.{ �C?EA  ��N����z_��[1ǻ�u$`�6]�h=ž�����H^1zח���a�+��O�Y��v�&�n#2�J�n �Xir���Hb��mԋYy	wrf�~�E�%�.��g���o�~D��U1�sn���{<_w|��k.��� v@�6�_������)'&r{%b� �'�3�͌ �U�HҖ��#�y�ƭ������y��RƫÑ�,U��QP�'Ѐ�&;oG/�|�#u�ⲐG��������<�=�]�Oc/8��4A�������>	��ʐ�<ý��-�]�E_ޭe �V���<	�o�N(�0ۍZ�rf���
�t&q�*l�{�N��D��ƶ��ڵ�����Gh�z 5������)���?�O5<�hV�����(��ទJ��|+b�"��"����b������y�,�o�iJ�����3m\|���m��h+��_��q[������M(:�fq�?2��j�%I���6gqs�rW�q�_�:�q9�j�C1�+t�K��L�x��-v��/i,�/�XRr�PK��~Ф0O��k�\T��%D�fb$�X�'�}�})�_I�����y��ܷ%����F���G�3�������t��j8�>ı#�cPnB�^f-|�:�շ~ժQ��ːJ��ׂk��:�����up��TE}r�ef���ǌ���>�gGT�Q�*I��X�´Q:f���K���xV�����9��aT����)�83����D��P���C��*������.�RK';��ͮ��R�ƍ��R@=�_�v^�T�g.��6��K�e�,W=(ˢ��t7w3���g4�-l�Vع�U����IAe�[�H�t	ޘ;����堽����k/���A����?}�K��t��B��hi΄ﵳ!=l�����p(�Kaɘ���!�1�Vm�g�,U4{�5�6��(�z�M�2-����E����csy���e�[������R����EP�	���U瓧�l��3e��F���Ͻ��z��!1��`�7��bUj�^
� ���&�nkZM?�6d`&������z��*g{k��@�݃��q�6؀���H�;|g�y�X�1M}��J����)���=]�#��9��<N�[*".���X�B��w�9}]��O"e@B/esP.q��7�hA���v�V~O�A��L8����D�؅eqNI7���<�gi�$�\��b�$�ҴDh	h�s�a�L(Z�M�?������V�����b}���d�J��[���O ��������+��zx�q)����p~�=�������,�{���h���ǈY�v R7`�3ęţ������lW%�eF�Sl� �S�R@����d�E:�k��a��M�̟ ��77r�D0��y�i:? ��?�"Q8�n>��̙����g·*y����Fl~Kz�)_�S�jTK���Q�҉lO�7UJ`7bb�S�=���V#��VTd�U-���nN�G`5i��s����QU�0�:��t�-!���I�E��0���!DE����w��V�M���LkL �PO5��A��>��Y[���,�����9��
H�l�A�_�>��L�nF
�������%�&)@:��kH2F�˻G��!j1nr%�S�0ǀ�os�5W�N�i
F��p~P@��XO4̖�)��@� �K�4b����ZJ�S���F"�)�U����Z���g˟Of�m�o�G��V�n"N;m�4"ks�ΣV|�C�V2oC?�t�����A� �I6I���
��|>�.!���`����q��7�3I�S�{�I�V�Ҟ�#a��$h��օl�CZ���FZ��0��#�~��#r0'���uJ94�6�� =9>#>i0�y�U-D�3��!Rt����k�it�k-����"D���P�w_:XU������M�y�g]q;���#�D�����%0ܚB-)R��h���堂r~��e��%k�v2��U��>����u��|W�=n?�X\�ϻԋ�[B�6�>	q�#4�P�2oS����9cp����X�|ݵ�ܜ�I�e����hC���۽�#S*��}��Ϭ����eb�e9&:*iJw7�&6�Ot?�h����i�T��W���y��#q�LӻPm�p?&n�D�t�u��Ѝ��/���| L��[���C�<�%bO���S*��^p��<�j;����Y��D����������&��q 5Wy������hkxf��E�Ѳ ؂�[���< �x�%6�V	񎜢Z�T�;�F_�v�s�S�ݟ!�c��%O�j
(��RZ �׿v�lB^�������+ۓ���:����ʑ8��@���2B�F���Y���F�E�%�Ҳ�S�o�"V��E�z�S��r�E[M9�\ۿl`20�d�. _n�?�Th
�	|�5[/��nԭ�q(l؁�5!�v*�wh��������2�Y�X��۝��6��5$����վɱ_P������\�S'�n�׬�s8B��[=�V�ɢ��X a������Ӫ�O|�]�q������gv.�PT��U.%c��&�:d�V�&����;�v3/[�r���힧�w��S�q�9���H��$� ��V���������"�b9�%�ˤP*d;GQ��A��bxv�o�k�nT��wm��mX*�����L�<�-��tC��8�����wBϷ|���Ͳ�Q�Q���H��c_)�y9�.����ڈX?rQZ�ݖ�c�#��{� �q+p~,XJ�vi��U�{�i��hO8��T�l+	06�1��}�zL<��Q��\F_=�8a`�]����R!4) .��H�sǷ��'<ʲ~��g{��ȼ�|�`�\ڒ�oQ���w�R6C�l��l��g��+ݥ��Y1c�[p/<Q�X�NzRP4���f~�Oo]!�F�w��Q����j����5��
M0�)`ݔ>F*��+v�X��$w�-�2��Aif0���h ]v�^#��c�m���!M�p8Ň��2�:֑�j��V۷�<m�7�2]�?_��>�`vG���{�4�r�_�8Q૟L`T�@u�=IG�l�L1Z"���3��q"!&�F���)T�h�����*���O��s��L�!Uc�f�*����r顯�Rz��îMP�=K�4y�2_�kѩ�A����>+rMj�}��ՖD�T4��5;-�P��Օ���$sb	�Cgs�9��wE|��˦H��qn0��yb�A����t�������x��ƕ�Nz�'$�z�@@ �Љc�J�&弹t�a�h\Nܭ�-�=�Yw,��z%V��1[�?����c�rd[�����B�(B�,G�7pщ� \c=���z��ܓtN�=�4~�"�p��c��q�?�a���l�S����=d"Dg���IÑA�'|�4,/�´�RC{��$���E�������݇i��I��?��^��}($a�cɈ�ζ��l��}~�ߚ��Q�6�^Ó��Br�S���̑�l~�82cw�q��'n����H��yF�Y�.��PF��-��Z����m���P�>!���)j�$ɋg,2@�)ć�d��j�)w�gv�`���� ���2��ԗ�dfD�*���O��u���s�1c%�d&��P���Y.8�ܚv�xmu1�y��P�����3��G�|Y�t�å�+��x�^��3o}�48�
�W��W.`��,��%@0F��i�3�c��һ�,L�D#��ǐFN�!@Omeٍ�ao�10+��Vg{كZ"v��f��ߜ�ޞ�a�LrhU@Ě�w��bh�-�:KI���dO�	�J8p쪞o9d�)xQ����K � �����7���=e��N/k���-|��d-�Rғ���j��X���NP�N;ё3�U�`
1�&1��$,I_��a� ������۬[��u=8�};H�M"{���:�����7�����uO%�:A,�G��9F��OW$"�#o�|g�[�C�f�r�\���}KnOԮ�Ta�*���M�A�~)�8.����\���旮��Gͥﴶ�
)ԺR)p��nxw��4z��;�ԑ��Զ�9��hȸ�����6KO،�?0��c�
�U3qvl�����Ǩ�:�5����D�?/�jZ=�K�E���m����Я[���7��h͟8bסj�:��|��>��<�;��·�fI���n	�tH�䌑&��R����^s�i:<
V��5���vw�,�>�����Վ�fO�������Y5��C<02 ���L'�����,Y4Ɵ�Ǹ�������J�]����#cZ�g$��(�Js��W8j�V��_a������R�w�$���M��lAd��QI:_��d+����&����9	:
��Yl�Q����������ƶkD'r?�9ФM~ڛ��=����> �n0ƺ�i�ҙ�G;���xW ��I���1Y� �weo(6$�
q�A�h.b� �Q�E��ѲL��I�z�7�[X���|+����/"<(ǀ�H|��z������h-�+�<� ���2�����̱��G%�X��L���b�Ң�R�(y�b4f߆E��.���V������<�=s5���IG�{�Vv|�I.ޅ���o@�)_�҈�/�)��{��� ?c~�z��:��U����xZ�@խT�mF��yo�u�i�ø��U�~8L'�o�&�6V/b9��b����G9G���T����<p�]Z�v/�|4����
a���V�	Up�wT�<�Z��=��I���W���w��2�{	�E NX!�T�ZV_��\p�����qkW{�6=��1�ǭDf� ��q��-!�h�c5�G��"ݽ��V�6�3�/x�1۝��g�2�J���+�z��=��S�n򸎦M����	#�JE������\�n�T���/�������6��=z�(a��q��$2����1/�Iir�6��{xn���_�5�q@d¶QIC䙶�Ҫ�Kf+�L�8�t��:�p�J/��XǇ�&�Kc��$z��˄\{�%"��fIs�X�S�}}"-ꈘ�I~ ��e��|�%�V꼌 ��J���uw�tW<���ϲ y���ĸ�{c7�m_8�-#�(��<h�-hQ�4�q,��U���n�I���m?~�S}ٗfD�uǳ>5�E�r���&*��w��'G���4f��K�H�x]���r.�� #�a��I��V�8���=+�C����m��C3�^4��9�R��/���p��y�r��5�R'M�_m�^��g�p��U�,�3���,^�wˉ��t�Zl�� g��.l+y���Ĭ��7�Al\��FtИ����2�W�?^�/�%A�]�&r%Sݙ�\K���6��%�H�ຒe�|��(X��?��R���bEmܷ,|1)�<�%6���(���MfkS����i�܂�WGc��:��׻�5/ǔ��ƓB��G��P$�ς���G�s��3LsW������Dnh��n!x6`��c�i<�j�&e��m5�ƃ�n�"M�U�6�0-���۩�x{���{2G��E�"e��Uf06�h		vH�P�g�5��1��僓��a_�C��$��]�O#� ���M�v��?"�s������꼭�*�m]�P"L�J/,�m.�7Y�)�bm�҂<O3:����2�~Z�D��~e?a7>��<@�k
�B��ו�қ��D/�#�;����D��3S��Џ�<>��|V�x�ぶ"b$[�����K ֞���9���g���4R�V�n�?V�D�Ip�u=�!��<49��5���l7v�5�N���R~?V3+�&Ū�#����3������d� ]�RNv���d�fO!��|c���/@���q�������;0�+y�~:&|G�xbQ�թ>%��3�w��?g��Cy�
�-��KA�e���S%(T���7���v�sx*7<[�`���e�Sf���3<��
�d���-���n5�o`�m������WwQ�!ͺ�G���?-(�d�0���e��p�c���/���9�t���Spk3O�[�5A4�3�� }Y�;�S���5�� 2�N퇹�}���!�n��#�g����C&]��p%2�@���+����n�j�S�3��"]�Iw��6i����\Z@�X���/̽$���������V�wf(Z�[��b��"�H|T��Z��Ng���fE��o-T��6�"����<�W4)cӵ��|�Y����Oo��xt����� YI��Q
�o�|��!�5>��J�ָ��7�4CI�BՎb�ue��yۼ#�p.$���̻ͻj�}��A�,0����%}p#���� u�߿4&�1�'�<>
�0k��UԵzº��!yB �ط�k���r�������WΉ�����tX��`���tj��nߑ;��C����*�U׃S@�!C)�gmh$/���9lre���,ء��:�v��BUN�>T�⟾�E��,1�$O�*�vB��q��R>Pʽ#[qoP�#o����~'9
��j�@�V��Nޜ�e����N�Jr:���*Sj���*�+�QӌR�e@�*P��7��6>��?@���*�J�W��$���
�L��m��(?�%sDX8Б�i�дu��R�گ XLč��P����3h����_�J7b�1 �^W�b�yj�|�j?����C6$��[�������� � �^"	�K�Xx��mE؋�Gۘ�bj��� ��%�.ƒ�0R�� Z�e�;����}��:\���	�b���U(	�ZGa��5�lI��Q������҇��F�/�'�O��8�����kBj��˘&YE�FL�%;���io7�&�B����S�İҾ*?[Ԩ�\B X�����s fI�?�J7h���	#z�[�5��KF1�#6 l�Μ5(�vׯhY0֍������Y\��"���]:�5+�����R�y��(�W�0�b�x'�Ή��̉s=9I7=OM PnUU��aSf4�%7���/�C�����=w�Y6�v�'��w}Z鋣�.r���ٖ:��í���Hf6vz�.[�����R<��}<�U�qWU��^w�H:�2��P�'~�]iJ���Ј������b�Л�2��*Ɖ�n�H��b_j�o��n�Epw�+O��<*���Q<�3��_�H��;�w�$�|���Ơh��Qu/rq�*/�)~q)����L�!��?@tSQas햎<�#����`�+��8,��T޽��|��p���7�8�\Y��S�+�Jc����}
S*<����FFS8(�]2����z)yK��w�s�ϸ�D�ʙ<��.�l�o��ߥĉ`D�ʒ��L��Y:,C�Y)췾*��߲����1�� pV�_3�z9������§�~p��]�h�F�>�x�����������
�(���m���&Fq"+��[X��w�9��y2A��1O�g����Ȏ�m���+�7���.
b2cvi�/�\#����m��<2D�?&�>T~pGoV��,�T�_���?B����T�b	ud>G�+L������C�B/!-���m�TI�D�va�汶��Tao�(�1!Tp!\O�b�r���Aj�)�D�K��5$ۺE�r#�'f�PyO���C]�@�LI�}�8T�7��PJ^��PgX`uT�c�>3�A�o^���\�[���S�č�)���dx�Uʪ��@%J�"CS[�{1'7%�?#�G���I��I�	���V����������N��-�u��J^��w��Grџ�������0"vG��u\U�H	^��]Ck9p/������0�Y*A����0g�-�����.i[�A���T�}�|`��YhJX�9��������v�����J(YLW���V�
�_����v����w�� $���]Wl�#�F�E_1�/d`�"�Ȉ;�Dv"9eG��e<l�����n�;ݴ�'Ƌ��'瀟9��~�������/�A�3�Ə)������\��]�� X��>��0i:�5�eD�C$7�,�V��.KN %CE�$����j~�=z{��[͹��jg��M��z�������EH��z���e�#�}�a+���u�����Ǌs���A��,X7����bB�ԧ��y�f�*�E#U�.����u��������gs��'�>�{Xgq|J��.��c�@��_�`Ȉ)�v{A�  t��O���^;U�Z}�I1���~�I�U�R�y����n�:�-�U��/�'���&�wA/��F��"��#�G�����v�%�<��q]O4�/T5,4�<������5�n	)��,�z<����ɓ-�a3��t�r����	��vNĆM۩��ZK����Zo�F�{�@�#"�bX����=��F��h"�v5����bB���d�����J&Փ�D���:}�J�J�+��ܸ�w11�Æ��3D�H͠>��J�H�fRW\���	Mv����ᗍ�,�C'��6(��cq֍�2��-���I^ۿ6�m�P�$��b�_0�qU����)C9�*��8�K�w�LGԌ�I�R㌺��2#/�W�Xno����K�t��@h ����\�A�%7�f��wX䀜}r�$�o�IA'N��5�>G%*�L�q���
����rn�	��,�y��M��e=��=�c��-�o�-�s�6�����KT�5T-��в-!$��nɤA���(�6N�~D;�߶ c��6-���/�B���ˑ��̭�Q~�;�c��[AB�3A ���yb����
�P'�m1�vnȥ�c��$2A����8�j���ɧ>D2�9�E�� �Wj/Bw�8Nv� �� j2�`֗ϚD$غ������׭ދ��~���������݈Y��z�Wی�q1��+�����V��GG���Y�뵞߾k+/���z�W3Q%4T����0��s���Ha��^9@�^;�6��3,�͸�u|��R�D?�qc�wN��u@�C\e�����E���mZ^��Bަ�k��R�q����4�\��@Y�y�%R�d�_� P^��g�.��\e0�hy�q,�t�r�teڮ����g�yl2ֹ۟^��o�A��^�&t7�#)Ӎ�^�P�&0'/�AbE�NT�J��bv��h����β����a1|�2x(��TɆ�y5��A�m�
,C�����'6E�+(�M�3���yp�)��3caA����p��օ�����aV�n��P+����v�}H�T3ӫ^�tL
��7\�k����!_�9`���$j���..n�Q,n�|M���6�����ϩG���?P@{�~�.&��I1�\�[6;����H/9Cg~3 ����1;W������#�*2c��K?]�����?吴���I�"܎\��>d��=���T]Dj�"��/�0._R7�)k�i����O��r������D��e_��7e"<̹�Rt��	�]~Z��"�D�b.�a��������m6�a���VBi���(bk����<�R�����'� ��l�`�h����o��_���k��p�=�u+�ž��z����&V^�uOw��Re��3�3��Q)ۊ��8����S�'�� ~ R5�;���d����e��@�;����x�����
d0�5[y[�:�_��m�:Q&��>L��:���jg�!�yb�c��9�K��c�@LSLi�T����])�zM��7�l�`e+[���S�
�:�l���d���-Tnn��8`c'w��pT�~��Qõ4�h���b~�-����X���Y��,���6�� �;dl���k�%C�5���P��Y�>����ᨍ������*�Z�c��(��nt���䝓��2&�a��׺�24�d��Vؼ���n�[�S�,��7�����|��i��ڻW@�_3}�ē	��Y`��n�W�bM|�V�Z�T��i��"���CԦ��ӬZR�?g���f���oT���k�"|[M�(�4�N��<��|�1�D�so�It"��̯ �} If]
g�|l�R!�*�?��톭֟�F7}uI=�9��ew�ۚ�'�#F�$�d�ֳv��1�U�����i0cx�l �# �\�'��ux��4����XU>��0�8NU���ى!��:��`nk��B����\?��PQ���O/�%p�X���G���;4�{;/�S�Q8�q�
ת����)���h�]��&�r�U�䓊ˉ:5vࢢUU�l>;dݟ�H��R���7ك�S�����֯���>7O?#"�!P�or�Ә�9Q[��<��+�������e����#N���M*;ඉ��c��S"�e��Z*׽�7�m6�V�?gMX�1Wj��W������r`L�Dm��?� kD_�Ǒ�ʀ�{�1���6~L+
k����e �����F1������^�%�.j)�d������*�b�����/��׌8� cp	���?�r�fxԐ/E����W�	�)&�j ��%$=G�����Z֢];�Z�$"���í�Ob,���.���(�tZ.�3����l�7dP�� �%�Dާm>Ҭ%i�6�%8|R�>%jB�)��2��Y�"�Fs�%B�Oo�`ׁ���ƀ��S��I���[�[�\I8���~�R'N 8�?vh:�	j;�[���Ru��
F�l�ۗ5�ziv�1�h���аF�=��Yc��	�j�$�5�YZ���:">n�:\��^@�I�*'��{ԅ�s�ń���=�pw��\	Va:[ݠ��黚��O���8��;F�d�Ӎ`��v�T�>���2%�.�(ĻTa:R`q�Ԑs�O�va��[�$�Z�l��sЁS�q� 6Å�%HAy�����Y`�z�s����Vb�;��9�<*�Z�58��*eb��o�%nB�Tw�����$*���}�<�j�Xr!���%����w��l|ɭ_n�)�Q������	�)ŘM������i�?�7Q?`�}`#$F6��t+��,�'�ޤ�|�C��8�|�89%��B)�+��]��<}���<���� �F�r�8�C_]y@� �)�\���Qs��{}5 � Bו��ֶ��̰�`K'0�Ї`���i� �kC{�]�����X��ߝ�8R1�a_ph����z�/_��p�	�|~� �]�F�+�?ݹM�����c�4
;�D������6�FX�++dK�XE��wV{ՠ`[AW�ēX�n_j�s|����m�n���8���x�u@�2�u=�6�a�C�wۥ�pmz�2˥�?��p>��G>���驋�;^,_���� ����T�YQu���G3COL�0�� ����L!�S��:+�T�	����>��Z��[�Y��`�ڈ!��fj���Ar�v�� x0��G�{�m���#��eߠ�~��*��$��i7�����M��me��D,b����-�A�����\	'b7[�C���v!��H���$��F9�K80�Jb����t;	J�M���������_��$Q��;@g-�o�J%�Ƽ���a⃽N�&4-:�.�y�w ��(E��<G[2US���3c��dɢ
s���1�(�G[I�p����WAc�ȗ�ZC���wt�K�=:��~dT�pXĕ��G�a�&ʚ+����=��p�̗��ejqB��v�=�b'/��� �{���$�\E�6n�1(iۗ���g�񾃀�X�$����v.䶫#0��m�~�D�߈<��D�69���� B`\�ˣ���?�~��ce�v�m�����v��y4.��k�PyD2��@�H֥��m�v6�lT#�
?�j�F���2n�G$C��jj=/w�v��2+l e��22c����D6V��d�<D���(�ߵ؄����~ϧ��Y�1�J���t���K��,��$�f��g�K�y<ҾK��ʤ�Sy�T���j��arǽ�7K�`Rӱ���S�a����^��d�]�-7�n	t�`Pl��_S���Q�o�Շ&�o��-|D'�1��w��DL� �؈� ���CH��̧��k�\0��5%+�>�yvY�kP�'���U�!��qc�'���x��:����n�<���5f�DkX&�0^��s�2����"�\�\@n��S�����ߟڰQ�i�]i��$�K��@ƊP�	(̑���Xֻ�w�O@��K�5Z%���6p="I��P���i��Z�n�g�hfZ�o��^�?"�]���4}\�Ӊ��|�����TLoft�G�9�� ��EI��
_'v|Y�f!�20l���S��}�7�{�I�c�6>/d+ݚMl�#<�$� h� ���>m��q;q~0�f����I#MX�����u��*4���{��>ކ50��U�nE�j�!M�\�,��k�!���n©�B�=�g�]K��RݎX��r�����HQ��P7;|=��>U�����N&�Ն�)퇿h�Y&�@��r9��􉠯lv��U"�W>�
*���s�������sh�JKm����Y��>��#/ĈPopgo�R˘��9�J�����2��P�����veaJ*�p�{���%�tI�*h�ȉ�?R�`p�`̈́e��I*$`�7�R6�?��'��W-���W�	vxn���!L�sm�NP?��D,1�Ј��O�ڃ��L0|�$�����`�ߦ����M�1,^+������j��W��-����N��&&������J P�z�27�󟔯x���E,`�:SͶ��sw� �܇%��{�1����N�ZCN�;�s��\��TA�<�1�6X�E��(݊�Z�]�	n�l�U���6���զX���>������T8��]���B>����YtDF��%�2/�]o��zF9��rZS��nҒ#�[(��\���ל�_40 ���?d�h'�	��[�\-�Xѭw��lӥ�5|�sv��h����]�w�j5Y0ML�v��1�75�W�hoH�˳"gSO�+B¶9�'����2��s�@;��y=#����0)cCa��u�����h���h��+��}�t���ڍ-��v���K�L�ߤ.����A��:�\y�{�\�v�V�[����h��^=\�n�q+Zò�HJ3�����ѝ�����E��u��y��b�����*b�B|���'b3Ro���n�rvw���鮁*B㏊�;<8 {ۥ�P��vB���w �|�`2��DژNQV�����~9�)R�v���iB�u�e?'Q��4�b��#�I+K��,�i!�z�PҴ��B�o38&�w���q+�aװl��}^�<�O�Wh�F��8|J�]�e�-��)M���-ȩs�*�*�{�m��ׂP-�C5M���`��=Z����ݤ�dC�MZ�-zl+�����m1�PGp*E���fz�0��|l��t�~�-I]���FA8R�L����� �T��PK�
ȉ��鸔yf�FŬ�+q��X��w��W�M$'A�
����;����<���Iml�Y��񖠋�����2�&�%_���۲�_m'�2��?z�@>(��Gk&�ȶPH���}_�2�P:�Z7�T�Hu8�G`�LLl*ٙQ����<�!� l�m�T����J�X��3�(+�|�w��v!��~f�+N����rd���-�v���P��Ú������%���K�n��h����,v�y4M�}����@Kg$|-o���v��)!Db�l�C^tՔ�+�2疧��9�|D�L��0Š4b�0���rt膌]8��:j��t�)TӴb66)�@ ���I8Jr�I��#�ao��N��S-[;(�|w�!��|}Ήt%[,��p�Uc�8�d��k|��e�(�+�G�sRp�w]Iac��'�k��w�t�;�=��m~�{2p�h��K�R�ua�,��뽫㨃=r<$�'��E�A�M�ޘCp����#/�F�ܭF�{��G$�0E!��c�+�1�iH�	�����k����v�$|Ǎ�?�غ�U�T~C[�ߕ ��j��6�T�î�B�~��Ђ���9�~�3cr�������n�c�y����	��PF��lJl�Ulk�L���#��Y+��ۅj�t���k2��$?�����j�OGw m�vu�Z_6� 2_<2�����cD�/�� ��)=1�=?a�����@��v�(cY�h���s�� 1�Vj���y;����G�X�Yp���~l�+�"@��L�3J�4s4$��9��RՕ��m;a@K�^�A3k?��ԉo���&Dz"B�NF�@)ëeT��<Vs1=�S�`�{���}R��!��߷	��@��h�=��6
��jI���<KO��.�d��%u���v9�yHxL���~U�ѝ���|�k%'eB��Nʵ����+�����[���6���3{o��>gNֆz3���`e�w����/\Iڀ�<f �� ���V߶ug�h�8Z��h�̀�a:��W�#��Җ@���[u�:��G߻F.�O2���^�R��g�%����Ʀ�\إQ}ƽ�O��T� ȡ�:��<_�)m�{l�\s\a2��ܤ��z�5ג��)���n3�z��.�z�4�i����)qg�c�M�2���� �je���o~�A�AEuU���a���>�( �P5s_��zu	j�JK���GN�Ft��v##��f��Cc�8�(�j]�e�||#$j�|$�WB��2�ڷ��c����	vX�H�;���մR��W�y�i��mV���5�a7���:� ���5@cLmI�>��kVy`lx혣�0p��O�#x�[���k//��r��y�s|@eEBi�m�Xx73��)��
��i@.�҈X��
dEU�
z#~�X�����K�Q����7����V��*�,G��M��C`$Yaq�sG�më�^W�� �M,Q-�y�ȾX��m.��\"������囹>�u��QZJ�FӏJ9�l�j� ��k4���̟�6$�H�ɁGW�P��Xn�%������s��K���8Q��pr©L�v�W:��$�y­�/=r+����~�ڇ��	j�G:�ek�N{�L~��Oݔ�k]�[=��_��_�j٬,���a��L"E甘_�9��_&��\��DO�k�abצ��3;z���;9}�<C���� ��D�` ;�9�H`G��K��;���,�?� ��L��K݇�Vb�H�c�m�9Y�;�F9�����:��������;y���f��
����p������d��S�S0��u8��T�4�����A�"�^U��i'ڊ�q'�OA�R�\�Ѷm��VC����hr����݆A�ڈ8�x��R����8#V���;�8fh�w�;Eذ��Q�̡���([������ ?^}RE���L��5Tb��7�B%\�3��
� �&9}��B�7O4X,N$3-W齩����
�MPoOhR��e�"��d��4�D^�W�I\��u�����~��1����_��dw�	gT����ՈБ����`�1��v���������܆�@���Zq��F���C������"����U�f��6]�E���>�7L�&0���=�I�~��	�kr6	S����êJ0������ޤ�*�@eB�r&���'h�NM3#���dbB�������?�GjP)�4�!Z��e�mMq�k�^�'=��~&�Y0��C�[������ki����wys՝~tf�Z&N��`p83�BW �	�F*!��s6F�jd�bѷ�!�'M�<��+�d9��RHZq�q���6��M(�a5��3s%��I'ܓU�Cl��kI?Co�s��WM4���U�Lm'�aB,��yZ�+�VB>��dc)4G��߆��6���u�`�e9G���6Q�:Ft ��XUR�Ԑ�>���������s�$j��t������U���ۇ%�`�38-������R�h��݇�#��'�z�BS�g1B-p4#��ʵՠPz�]��PƆ�@��x���;B�様Y�T	���蟜"s�i�ߏ�e�zh�]�= �pi�xF*����ADE�.(��m��PF�WRm>i��7���!;�9 �%E�CDp�����&5�^ '��Pe���`�CI���tD�iэTӽ�YN^n�!PSL�u�3��*�A�먪Џ����6�6?�Yr����6���/xP~P�x������C[L�-j�%V	9�3����n3I�kg�`��Ѭ,��)u{��G���Pu"6^� i���ыms	|٣�#�"�h)�a�,�yt�^�zDC�0�pr���Y���zX�0�����������-�w���x��w��L��JDcɩ3�k�̵�H�w���J�3WýV
01_�W-�~��t� w��6$�>��n��l�w썲ă_�'d�r���.��9
���3�dl�#],~�Z�	� ~��wh'S�69��<~���ǲ���R`h��{�3�����Hݦ��Z� D���������e0��$�A��B�s.��� )EI�h�͕C�#,zgǆ[9h�}���>�C�p�����4���H?z�HL���͌i"L+DF�a���~���vz�R&�Xq̳�׀b��{ԓ�&y��f�]�E��).��<���ܡ�g��]��sv���J�{D��|��K.����j�@��[_�M��{�)/T:{-Q� �Ӳ�;vӌ�U�{���Q����ݭ�L��	&y]�Z�Ùg�U��Ylm'��&C�z/�{��+U~�qtG����!���<�bc]��/@D4I)ǁ�xr��f7	a�ʘ�N<�jV�5!�Mnf�m��^���)	��rN0u�ەA�Z�Hv�݅�|�Ζ2��{�肨��������r��#,K�'�h�zY5��N������W���p�p�f|�0_��1J�t*+ji���ڂ�#���^�q��4�1�qJ���e�\�F��u몤p���g붗yϿ�������(B��q�:�2�re�I�p�6o����N�y�_�|�qA�<�r��C%�E�3zkK��L� ��5�����sq7�/���XZ_����zK��Ь`U����\\1%#�'fj+XМ�}ޓ��	6^I�˚��gʓ��%B���z��D��;�7������������Ĺ��cXr���-��1�"����Q�t=�R�a�߭s�����V��#� ��}z�fNǔku�FUN%[�$�* ճ`�[�Y�f�ԢK���x^�t�����A��a\f���K8;&����$h�������N����o�t\RS.��#�L՗��Z�W��Q�RH�_�8�^�"Dg'�����{�����,_�˪�pt?,e�g<��l�N���N>���}AmZ��t�C��I��=� �/��xA�̶�G���g�|��Jtp�Ό��)gc�r�����(��ɠ�ӓ̠9kWm��
,]���=ز6�<(�O	MǨ+��f
������c{��� ���"7R��A_��P��ȕ=Pū����9�ie�t��3mg�N������9�Ԃ�d!9��`Áשj��j�Jb�ׁ'4�ns߾MG�6l��՛e���D�ٞ�{s�h�H�����C6���R�H�ևg|��`%�1U.��p<������ �]�FP�A�a��A��c�]"6ށ`>�0r���]�{ "mL/m �.y�M7�W����'�Ow2��G��S�D��-ey�7�
�<����,ۗ�#	��Ҽ7FDp�8�{�E�T'ƵU� �G���w�7�VܓE��5�b����l9)���X�����*,�Ɠw�����'��yw����p��M=���������~���p����5�&�NR?�3^fū�]�'��t�mw`�[�E �S�RA����d��3Bx&�����U�H�(���?���=0�Smy���:Gl��Gl�Q@RT>���ԩ��
�gֹ�y�kʾN@K�p��1U"S�!CTS��ה�뺌�tJT7]mS`??���S�|���v��w@d�E�-� DnV��`=u��y����JQ]m�B?��|��-)���QMV����ѯM���6n���`U�i�T�lkTu��5�Ů�Fn	Yc]��4���ТA���o�tVH�gK��nNK�������&1D����2N�s�Okż)2{nz�S�����̟'���Vdi��x��@���WRS̞q3���w��y�<����;�ZRݽ�\�"��]�ٕ�;Z�x�gӼ�f�+vo���^�R"V�݇��4*.�����|��J�^c�oKF�t�l���*� �S�I���
�+ |F1!~L�g�� /e�y9�7��I��T��?�QV����#i��$p�֍e��Kt:�$Ob|�0�.�цg�#z�u��(uR��4ٞ�( P>+�\0�>U5q�;��!Z����k����s�Z����*������X];��!��U?�oP�;�2��+�Y�T��]�ܢZ�)ZգhU����r����m>�-iKv:�~U�0�>u��t�����E� �`A��A��=�&^�>�q#<9�P�
o?ј�F�9k~�����`}lݽO��e��������½�*� ���0��!�m��eA��*qFg7�:6�mS?�G��˜��\��W���%�2�+��L��Pm'9q?.��D��6�}��Е�M����ЈWLt���KԬ�-2�� �9�u2Y^x�t��Q�jCb��а�LKӦ,h��	f��c��&� =�ڡ��A��g�xn��E��+(��cE��N ۝�%>�{�^���CZ��y;�й�~[�[(�)Z.��so�r4(���Z�����lJ��������&�3���N笿���C�8�y>����B��f�KbY�	�F�d�%����T^o E1�'\��>)S�'��q[U��\�Gkh���l�� gY�?�Z�hר	��[^z��~���Tl�Z5)V�v2xzh���������Y����6:�>p�5,����19ю%X=M�ː�=5�#t'�U��/�s@ <�.�=�\��i� �aFc��A��S�����q�
��������Ov�8�X����K.-W��.c�:l�t�.q����v;�~[�LT�������[��q�����E0H�^1�`#�I�^�����ɒ)�ITbA����l�*�-�O;��I�b��o�x�n\j�w%�Z����*�������<巵��℉�	���KwJ��|��Cɇ���K�Q�P,X�k-�)�7� ZT��rU����?!�Qb^;����#��V�(��+x#�,`�b�~R��]�n�q-8���\�e+�H�9�X}��><�9���Fgq�8i$]���Z8I)撚As��oׂ�ʺ:>�o���К��&�`��풪����bk�Z�C����1���R�3����1k�p7f��`S�zZ�����#T�~���]���F���Y{���]���o�=�z
U�A�1�L�F��F2�+~=�X��w�[`�: BAqd���i�G�f���%<m��)��x�ŏ)�2䁢�Вh�Qۿ�{m��!2ezR?g�g>�n�G�kȃ;�#�_���@dG����T���u�ӿG���L9�����.��˄!.q����T������2�������4�/�!]��f�x��Tr�Ga�Zl`��Tv�U_l����<���:k���z��o����[�F��Mr��"��՞w�\���J-����N��|�bBC �{�A|#�a��η��	��ym0�yGb�"b� ޞt��@��ϼ'˛��+�/ ��ǧ��fz0&6�"��Wd9�i���W;�d�7ʻCj7D��z�V+��8����'k~P7�!��hC�O�����;ǋT�z��^ ��P%�RuҜ��|]@A����7ԋڈcE ������$>x���`x�冪J���j�`��[�ڑ�\�%hV���-�GH�I�wȈr@M��t˒�qBG ��*�8��qu��s^~޹�,������@@�Yz"��S�����2E^��C��pmF���.�24�C�?�̶$��gq�-�sw[�$����m�,��3�)���J��N��S���$��6�>.i��Q�J�32�U�N��?2�f��k:�T��̲��=�����M���TX�j�%���䥿)���7�5�;�i����r�a��H�:Ҏ��Ő����r��l;��~�[�|m��y|:
/7�TmLD>��3�&��gصa�퇱�ь������.ar+�"�����A�9���&�W����]!O���a�`c���3�B��g';�n�<ɫ@�	���Jz� �"���H����Q;�h���ڄ�fW�L�'�R�V��H�~m�VV�P�9�$G�E���$F�76�K���"Ul���l�ݰ�p~){�e�:~��S���������'�[��A66��d��/$u�"��_��X�R���nm@��V��(���DɆTcB$� �r�-?���GdV�;� %h�@���&i�-%dQ�'񣩗A(��l�aLд�O}t�
T��{L��8
B�}��}
)-��,/�}�4BVe�Oz6QN*��W�E�|Xp
1ߦoU"{_������d�n^�J�4W���\B_���mQ���1]k��>�d���	mG��i[C��$�$e��fc1���v%Bj0�x��'�@_ƱO��aq���Ћp�kV�%J���pع�8�]�nZ���޷&��[k=�.ĪD-	@��r|�S��尙>��,
�A���iI���L@��rl�����Ƅ�e#�̪����<���P�Ę�V#�PY0���Z0>N�T{Aq�Bi^{�W=M��&0n��9�!��Wy�k�����s���t�u&��R�8��W�-���!��|s��F��fŨ^�'�MS3D���Ҁ��]�����q6�%�?A���~M� ��{�y�'��èɴH�Ŋ?���9���)�4ʋ�U�a�'w�,_c�y����~�g����4\����A���j��5��^�����( F���Ӟ�tR�5��]܂u���Bs옎���'�L��c����ݿ�M�`�-�����W�����i*W��4zG��ٜm�BsGA#��r��a�z�� [Y������,#"�B3�৞��T��R��#�Yw�o�a��Ĕ��Lᣅ� ��i��*T���AJ�7.��������WX�i|���;����+�C��sD����V��,��$Y�'R�P����K�CBY���y��&|T�vN'^�~P�ԍu��@���Asօ���Ί��[5��/��7R��m��TGix֎�����U��.][��xY�j%\����(S�;��Is��f�o�r;��(�����ʦ�O4Fu���^��� )�Q�������C2"��'�ج���^N*C�llp�.��u�;�b�Y��T�@0Ym���>	����Z�Fd��8d��RH�J
yl��nq*lu�NN+�F��J��W���VK�_V�T����rw�&�$J-H����l�/����_��dR���]���a9�Nv���Hl��c�� &Lݦ�Fƽ��'YN�9��I~� t7���v�*�Ή��"�������O�" �DK��2���m�'Y&ev��$�"�#9.	�e HyMEO����[p�2z��c[?}��C���ā̿��"������pdH���z%2�����/u�+��ԧ[��8��<�v��$GN��Xw����9b4�z�ه�y��fb	�E
�.�r��/�L�!��Js�of�;�{
��|<6�.�t]�n@�fX_�ۈ!J)5�{��M fD�́���!��U�f�;�%�ǳ���r��y��<⠆�ß��U�"$�ՠ'��&I�./��ְ��� ��G �T􄦺��K�<��]���/�4������	�}(��@<�~�;PQ�~A��疤ٟ�k�	rE<N�P��ۍ-Z�U����Ͷ�x�{��0���T���(�|�)��tzhϲ5����	����S��� ��Q������W�,��J@�+p����iqʏ��ގ8-��_�0��JL���?1\Ja��^���d��mX��?�.�5��DO%(HEq���2y�\��/IЃ765$�B(���_���qn(���.Ck1��93K��L93��{���+7�e/ߋX������KfOq�2������\bw�%鉤f�#>X.}������I3*��ז���
%���c��<���Ac[����d�� ?1�Ec��}�+-����-GH%Q�o��XA�٥�v�CDQ�C���F�ƛ�} �8fK/,ǚu���4����j��*&��&�U��f�#K�v�x$yD�rI���Mab���Lr8�B�D��*�Ѝ����r>���O�]8R8
���+�`�l���5R���_���^��g�0�|;3v����,%��0,t�ؘ�F�g�plR�x���Z��A&A3��~fatW��I��Ȅ��.��F^�/��A�{o��HWڈ��xM����0��#z�/�����\�#Lc(���ɦ/
��{��k�m
�,c r�S�6e(%�,M�u���Ul��l�Μ�c�����zy��0��l���ðώi�PK����x_��F�:
�3�%�ܔ
����ϋs��B�!�~`ɭɩ0��j(���N��-�Fn9�M�:�6��Η�m��g���_
�{�|��N���i��|�?6&I[�ʼHOOg����s1[9����K.���J`|�>~]�%��9������i�q"��g��H����g�]d�	"�):/��E.9m7��급�D��hO���*��%W�DbPee7��0</>�r��)%���Ba�D� ��tN�+��b����`�#Ӆ��kVb���v�b���2���rf���̓ �{��p�ψVv��M�f	닭ap��=�cM�#�o���<�Z���$�v 1��U���R��M3	�q?U������m�s���!'� 8h�RU海kd����_g�)�[�a��Ĥ��T��X�0�G{y{m�:�y��*KQF٨>l(�Z
E�{�g�STy�F
��sKK���7��Sl��T�9����̍:�7��4`�ɣW%S����Z#j��td�+�-t�|n�`������weQ�?���b����-�����1tZ����ΈV/��@�[M��k���c_5��G�Vd̌�Y�L��:���ȣ���y(�)c�z���-��H��n� ������&�[˳���2T���%����n��@S�>N�W?ܟ���Ȝ��i���>�@�!��̤;��y�*֎�Ȃ�y�ޘ�Z�义�"���c&h��i�Zr�gw$f�.)ot*%����"�	Y�#�r4���\w�|2���d�o�tBo���}| ��I�3�
2�|��4!��_���W)ֿr*7�'�I]�ю	;���I����#/L�$�.=�ӄ�Q|���,�蝨0$��ь�#@�v�G�Hu�� 4����U>��0�v4U;��� �!��q�߮�k��d�9U-�|Y��p����qM�E��X���g���[9֜5�c;O�J�q�y���ʊ �(A
)��h�����tr��(։3��v I�Uu=�>[J�����r�W�˱@���5��������>W#B%P��No�D����9q�)��"���1��2���eԐ˦CF�ч2��{*[潉&���2q��s��e��*���78�h6�8�?�s��QA
��}W�2�:K��l(L!)m-��?�f�D�?���Л�Q���V&.LKh�����#��"�f�M�	��r^�_��%��jI�.n��a<�J��n�O4׬�� ����;��+�x���E��.P��)|F^� !�*%D�v�$��g$Z�p�;��}�D�f��]>�o@О�"N�8��(0FZN�ٿJl��
��@�U�9��D��E3;�V�g8��Ձ^;hBx�R��Y�F��b%b�0�oS���*1Ơ�NS���%��[�h\iB��Y�r9r -�?7(�hZU�	�]�[���r�U�*��l�<5��v�kh�Y������]w�Y�7��)N]�Dp5��(�;K?��^�?Z�~��iqY'��ԥ�Es�?n�^=������|��aZ)h�)���p�;��ʇ���f�����k�v�[�^���Rb.�❻t_ :r"������o�Wv��}[��(�z��1��Сq�q��åѢHac���g��ܝ$�Cޚн�[��b���Y�6*ͨ�Uݝ��b 5o.'�nb�uw�3�<*�L$��H�<��5�x�[��a�����w�F|"c�����{uQ���ug����)����}T�Z�(r?'Y�Q(���5�
#D0�.a�+>�H,�f��eh�c{m�7����8Y��bˮ+׮����!}�$<�[7���F�, 8�AQ]��q� �r)�&:�� Usՙ�K`�@b׵�k���Z��֏`k��� ��/� �C��h�>*]��
��%��8B�1���p=z�&�z�IR��Ƒ)��~��D]2KF����_5��mX�'ø��N�
[�������̀$Fx�+���Xet�wv������AwW'�x�=����!m��+�m��B�� ����Sŕ��2�;��V�=�cV���Wm��r2�?�?�c�>��G^�%�	T��[L�_�4��C�-�8TX$u˸�GSI�L���\���S!�i��Z�T�'$��~������{t��/*���!#��f���2ތr�x�� �C�"�î�:k����t����2b��F����?�̫+M�Kg(���d�o�Kl>?!-�A��*8�|S�bW��C&qy�Ӛ-�������?�0vb7��&t[��0-�m���V-�����mȫ�@.���1E
JEH[���a&�N��-Zv��gw ��H;�\![RS��gc��/d�l7/�P�Y(�?G{#�p���9�c�w�z-n�3�t>�=Z&�~�N[p-��޸��8a1�ʺyj���=�C/����ԇ���5���ʂ��/��� �{�	j$-d�E�F�V��|�i�%k�ιE��Ӳ��>$�}@ɖ�H��� ��ׯ~��ߨ������6�����M�B������N��1~2��c��_������dؖ`�yT�?��QeP�����h�����l��،R��*�j�L����2��n7�K�24�j��w3/v�YRQm ��2>`F��
DV�)��Ќ\�ĭ�*]��-����ўgߥ�Y���j�$����1�^�]X��f8��kG�8hY�Ú�Q��+�m%�l�H3=�>4Ɩ%���ey�zKb@�!@~�)�(�e3^fF�'��z�CD1�,���   �   ލp�F˸�$�R=�1�#l����O�ToڬrN�'|W�DC�O���]�e�����:Vؽ�Da�w5,Qlڿ�M�F�ilZ���T/f�l����!��TI\&�L	���I!����һi7&�����o�x��f��T8���,O���bM�HR��V��x�Il���>yUJ^2_�Y�C�b|ެTf!m�04Jܴ�M���F}�*�K�	_�ts�\`�D97K�p��T��B�	5?��0�)Ҿ����6`�C�I�m�̵9��]�c�B�L���C䉹|�z���#CR����_8D��C����$h��ѻZ�\�)�Y E�C�I0<ĆDY�*]0�|9�)ˀm�2B�	�V� 4C�l��,ŌD3��!��B�IY �z�ꊘT�\h!���1ݰB�ɯ>�h$3�Ꚋ7��H��ZLB�I���I(�JX�t����`���C�ɖI��D`�YU��=��@ax���>	$EJ�AF�s��ʻN���QD����O4��V�d�27M>}b�ǚ�ug�O�� �J�-D�.ez�,/2�\�@��d��O��L�\�4ᐛ,5�șv薹���AC�>Q�1�S�#<Q4��-}���"��990m�g�<QP�I 2  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   5    މ04�̐��%�R(O5f��p��'l����I�l���   ��@ӌC�A+,ɘ�I'\	~�`%Ϲ>   �   ލp�F˸�$�B��>�1�#l����
�޴Y�:��O��d�����	�����"fŰu�pph��^�wS,�ش>G�6$}�8����
x��ј�R&?&����[���x`&�j�"<�C~�����Y,~(��v��e��W���%���36ڱ�-)?aQ�E��7Xp}BJ�8���D�5{>���N�!��X�Ӻi]�V�Ϟ������ē��.�-!�ph���Ȯ.��x�ȓ�V@".V�>��`���G@�ȓ]d|z�	�i.j�i$e��N9�ȓQ��
��p�GCO�kk�����ZG�<��"��(VX��N½,�V=�eH�<! ��/q��̂0�� n��iI@�<�P��i��`���?��%b���P�<��*�=E�2�:C�"�D@�0b�M�<���c�P�Cc٧o58L�1%Np�<I�"ϧ3��m��->n�a!��o�<���f���'$«h#�+WfD��h�'��Ň �¸��O�=y\������I"Qf�n�󦹤O��7����rX$��N�1^n��6bD�_��➀��I0��B �3b�F�d���
q�9�'t�Ex�}�'�R�j���2������6�|���'�L�k@ ��<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&�   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ����Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�   �  �  �    B$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�U曞@�VM�P������@��P_`���'4r�'d�|J?��f�s^hy�&A�x������ b�8�`XTv�|2���,�
�*��ڹz7"a��iRȖ:[�Fi��	�[ڀ3�F�\l����S�
��0ɂ��O��d�O:�d�<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&��|�����$��::�i�V�%C���e�Ԋ!�lK��O4�$�O��d9��~r"&F�L����� �45`� ��A%h�d��o�&=���1���Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�Y�P�{ � T�>�@� D�(1! " ��Eɵk��<�s�j �M{��$�~��A�(���4 ��7�*��2��y>���=���O>˓ I��"��ߣo��u�)9?Ԡ��F��r����y � ыU6��ȓ~�p�k%��^��1� �
$F��ȓN�� ��啦 jN=H�Aއl�І������(����� #zy�q��K!�2�"MF�����X���KV�w<�%2�M_�I��$�OD���B<�����J��`9���)�!���r�¹�P�D*/���2!�ah!���#S_l$�f��dQ�ݒ��߂*L!��F
�L w	�zE���'�@�H�x��#���P�P��Sap��M:L-���J`eEx�O`��'=�)� (仃'یBx��"���6�˰"O�q@�	��@�aKb�1h�Lm�"OaP����`��\���3��"O���lr��-�3|�z)�u"O��vJS�-��H+A��usp	A��>i��)��1j�L�B��ΥjՈ��1��+���'*T��d�'7B�|J~�A��99�p��G�fp�3�C
Q�<Y@��d�f�B;R�&D�S"ML�<�#ۼ|����#��(���H�<)�MםB���5
�=bxD����G�<1�Ç�;i��aڡb`�Ց��^ܓO���u(�O�=�S¤�BHC�e �s�۟�&��)�gy"lG",*Ȼfc�7hs����)���y�Q^�H��0��#�$��y��O��z�1�
��} ���qAϬ�y(RC��U�?A���I2F��Pxb�)�Ql��\�pH�Ĩґ+��F}Ҁ�:�h��=a0�A>�R��g�*� �ȝӟp�	lX����O�N����ql �Y�b@��;D��SvA�zb2��Kߺ�
T��=D� 9`�_�#X=R�H�8����'j8D�8���_���K��X�Y�(�RT�5O�DyR�G:nJ9XC�+����W�L��~2'��O�)�Oj���>i#�\��:�b��Ǒ8���k6`�V�<�fM�iH��&k�T5P�Gi�<y��
i���uA�&/<�� �Qy�<)��8
;�9$N�Y½�eQZ�<�O�3��2&
�ڵ��QP���k���O$�9j`&15ʱp%a�m����I�h��������v�)�i	0�
�ː���3^�M��LGk+!��;m&yBQ͓�`���k��H!�d�,PD
���/�|��Aɂv%!�$
ZO�9eD�J�΍�s
B�!�$PGS.]*��;��xH�jqO��D~2o�:�?)�O	�s�  ��ڙpmr���[��R�|�����I8)a�<�7.G3@O�t[�/�Y�C�P�2��¨-��X�΅=g�B�I�x��u��
�&%^��#�
�T�vB��*H��!(9�`"E�^�hB�ɛ0��!�@��� h�BD�H2�Q�'7�-A���L"<�X�a!���C���&3���I֟P����#��� ���9�h��(�+T�B�I�-m^��qJ\�{戔s�/	�ZB�ɸT]&� �Q��\�Ї��LUXB䉌v�>���Ã6Lh8��l�p�J��D�q�'���c��ƙ��%P!�ۢ��(q�'�0�K��4�����O��[�$%h����$u��	��[�$`���&�A� � Gt�$5.]�t?F�ȓ|�@9�e�-Dy���L$A�bф�b+����`�����lr�ȓp��$0�&��i�w�>�ܴ�O� Dz��4&ɖyy�p����>'˸@
�����	��š�O��$+����m�����.��"��b�L�yRD-k:i�4O�.0E(%l��y��X���놆�
}\yQD'˒�y�g�m}�p䃏�z.*)�����y���==u��AK&q��ih GȊ��'*�#?�E����ܓ�L�hFa��]8��!�=�?AL>)�S���'(���Z#��hi,���f��MG!�	:��ѡp�Ĵ3&|���R*!�$D(7�习���@Jm:�A�Vv!�d��>�p�$ =J��9���+#�𤜠
�\+%�3y��D�G���m?\����
=��>q���^ j�`�v�Z{ج)!���?q��>� �8�G�?��L[�"�)b��""O,����s�����E�<��"O���QfFI�Ѝ��:{*�Z"O|��ä:/pCs��~����'B�<�ޯW5� S���2.�H3L�{?Q��Fe�����'N2]��`d\M�֨H�@�!qg����:D�(�GزV����j�+��E� �#D������;%���s�f�$.A�\I®!D�TK�b�+0���딡!v(I"�>D���hB��(��EƬ8�<�!u� }"�4�S��L�����J�/vJY[3D͜<�q�OiIAI�O���3������8���Y��Y� ��������y��E���[�G��jP��!Ð��y"/��x�P)X�e�H�R!�Q�yJ^��qႨ��a �1бnD,�yBeܜyd�� ��*� ��@�C��'�*#?� �Ꟑ�g�J
�pt�2��4�>l�V��?!H>��S���DX�^�XCB�Q,�$2S�]�,�!��.�B��#$Z:a�*�w���W!�d��~�U
Cd�=H��e���v�!�DM�(������E,<�Vy�Cm�F��ā+M����G^
xL"6%".��$�>����X�s�, �W�W�}��5[����?9���>I��� ��p�j�.c~��R�cGS�<��C<o�y ��w`R�+�J�<.�Qھ�Jć!�b!�*E�<�2 �gm~�`Fĝ`��;#d�\8�H����-�L�ە��> �ݡ�m�F���I����\��Y}��Y�5�آ����9��9{����yH��E(
%Q����4-�Ա��yB���J�`��)�$4RJI	����yB�[�g�X2'm&t�H8�hO;�y2�6Rzp��Ag�@بCoA:��I��HO�$�zwΚ�����$}}�=��>��֑�?y���S��q��yC��1S��Vi��C�	�N�NhT�X9T30��Q�ˣ8�bC�ɆP�ɩ�X�"`n�(�+�%tB�I���B�aҀ`
t��E�I�"B�et@�@#� ����G�U��X���<I�� cNxԙ�	J���:U�C�4���%���O>���M1��%?|8�a4�������E����s�Iy�G5�&m��[�>1�5C�D�Xu�QF�"��ȓJ8���J}R8�3D˺%����~��m�5L[�\��`6���҂�#�#<J8G���
,�(���:F�x��Rɨ�$�O0��:r=��@�շ9��Q{�M�@�!��]1 ���q�+�9`E>컕k�NK!�Ev�iP&�%Բu�a@Gb,!�_�vpi�CV=��1�i�-%��xR1� ��M�pk��<M24⃋��\�X��$�"Fx�OL��'���9L�r�&��v84��H��$�C��$q��
Ѩ�9#fԨ�j@>1C��"h��E��/לA�����%J+�B�	Lb9�ÆȀ	#8t�V"�x��C�	�q�z0�e��#�|5oZ!P��'�"=�z����2cj�Ј7�ʕ�F$�R������OH��-��	V,MQb�ɍ�3�24A��5�y��٤#�4��#w�H�jA�Ҕ�yB%A`�V%�q�Зo*���
��yb*K$���΋�R����m���yr�B���\C��#K��$C5����'�l"?�rʟ�˳��8D~�� E�MF8��O��?	K>��S��򤗗g��AB�˾`{"(��Iս3�!��  1��e@u��8���H���@"OԌ�e�^�2��KE���+����"O�Q2+_�F	f� �H�#�ܤJ�
OV�k�3+��2@@��8��e�����O��H��S+�~ ���ͼHqh��v��!+Fȵ����?	�	<t!�̇�: �A ���E�4��ȓF��dՋİt���Õ���q�����$���7(ܣ�����'�
@����+O�UQ�*�Qo���r܎- � ��I�(OD)Q�*�)>��y�5�Y>}~����O�rb�i>}�I���'\���צ�1�P��-P}R���''�e�T�;n�z��Oչcb���'c����f>w�j	����X3�1�'x�`�􇎋@.��%�8f�t	�''4� �=/z�B�.�3W�>�N�h����)&U
n(z��N<3A��IK����|�����?AL>%?��S�T��bP��N��@���?D�$�f���T�b9ص́�?U4Aa��>D�hơ��b���'#˷Q��v>D�V٘ ��) E�s���	�Z��y��Y��r㨚(g/ tȱH���'��#?�0G�ן��$DٚR+��3�Y�&��D��?�M>��S���=4.� �偙�s�0%�r�X�E�!��<A��#wA�9��h3��be!�S�c�%�%Y�v� ԩؓG-!�d.]T��4�hr�`M$���Ȼ.������-7VP�1�D�_���䑞u��>	sg-��"�u�2��!���7똰�?)����>qV��
&�(l'��#iv�r�jc�<��aA S5Z�颥�\�>��q�_�<�aP� �n@�6��$����K[�<�C�x=\H�&�P��0jN{8����dF�q��)�7G�b*����L�/����n���ϟ(�IC}-'hpZ�
(!�[*C����yBg�0�,A��R8&�H����$�y2�Еf��͛���+"P>%�!�\��y2��:�ɥ��lr�@p�ۥ�y��Y�"�����m�+Ro�� ��3��	?�HO�2��4�S:\�ҁ�&$s�4:1�>�0�ϵ�?i����S��/�ё��~\ޠp��Rw��B䉝2�8d[0΄ifzR��bM�B�	�p��a���)C�j���k�Am�C�2i��5mޡoX�Q�gŏfKdB�	4%�]H&/��IDT( !D�hJ���r���E-/��8{���#vî*T�ç!ͤj1��d>��O>�|��������pL�Vc�=�y�ȓbTȁ��N����q���T�O��#*`88soK�F-|��g�1m�,�ȓ��e.؍\�nMb!B+=L�a�rt�G���;jd�!�V��e:�=��r�D�Td�]�8<	VX+8�*\��j�/XE4���O������t}�DÐ�:z��!���M�!�$D�g�����?q�8;�-g�!�d�U��i[ �F&�ƌ"�m߬b�!��ں�Kg\;� �6Ώz��x��"ʓ{j�P�S��)��a�D�5W���E��Fx�O�B�'��Ɉ8�
B0���!�dJ��g�JC�ɪ�AH��ep���GKǋG�.C�<7<D���>�Ȱ�7!B.Y��B�	�i*���M�Rf����şz��B�	RYРs��P�P�wiɸ ���'�^#=��얶g��m9T�X�	�.��@cQ�D�7� ���O��O�OW�s$��)b�����?&��'G�P�&�"���a��,A���3��� �]ytG[�7���V��To�i�v"O4P�P!M{�h`���h_���F"O6I��*�<6���냁�E^z�`��d]�'�fX"��V���R��T�l�%���Jb�vje�'��'���Y����,J�,�@���ܖ.X����*D�� �mδ��S�Z�65�'D�@c�b�*դ�%��Mʬ*p�#D�|���A�,s�$Zu��k�֙�'�+������v���IcN:9�T��m�3XQ�$�@F0ڧH��Y�)Z�Xl���J�J���'���'�~���$j��`9�c��z�0	�'aRX��e��$��Hi��F-Y��1R�'y�Y���%}�DI U�?_h|P	�'�f�
&��F.�]9T�P�Z6�9�
�Q�Q�{��s�u���"i2re&�i�'m�Y��h���O��V\�ؐ���%R�t�>o^c4c�-~(�k��OpTR��j�g≽[т�H��F�w�� ��@��Y�v+�6.�`j�'R&�A��4�3�$�_ Y�%F8�$)Zi\�|��	y~�jҸ�?ͧ�HOL0D*�a���8bH��Ft�4"O��vH��29�g&�\2����>���i>���_}b��h`�hrV@O �zH�m^�I���
������䟀'��O�\�("mV�{�DՒ��ז2��r�N����4OP�{[��X��'�d-P��ҽWh�a��s�h��Eʟa��]��8�J$�'��	��i��?ҙz&��
L�2�m���?	��hO�c��(6�l<�|��a[9��Bi9D��4 X;��sE\���Q��`9�	��M����'k�����-`d��BW��Dӧ�V4=���'1�'��Y��!�{Q@�Y�'�<l{BJ:D�h����355�����	WB([% ,D�(B���i*lAT����iiG�/D�������L�Y��T�&3ȕ���.�� rFD=�<���`��C��1���LdQ�(��#<ڧ%�M ���]�Dmz� ���1)A�'o��'�ڕ�P�H
�x4�n�@Й
�'P���j.X�F�B
�{�@���'�b�Z�m�O��m;�I��/����'�����t���� 8�(�Ǔ_Q�D ��!\<��d�m`���Sͮ���)��|����?y�O ���h�-eڴ����L�1&"O0��Ӥ� {v�q��øq)e(�"O� �2͛1���րQ�(�4x�"O@����$GM�[��[/u�|��"Ox��e߭lh�QP.G��p("U�>QT�)�S ��M�*�h�´���=����wb/}r���z��'ɧ�'>/�J� �7=~th�O*�,��zLi��L�j�x`�u�P3�D�ȓ�0��1eӘiA���g�?�\��_��*���K�����+r>1��M�BuҦ�"R<f��clм"6܍�=���I����$�<C�!�JE}��J��"VzBL�Id�I�"|�'���vDL@�pPq���Z���K�'|X�顬�.JM�)���E�R-����'��H�B�	 P*�B�K	�BY4��	�'FŃp��3L��m�$�B�:��
�'\@@��ӻ+6�Q	A�ۡI�0�q�{�'W��9�'_�2�����7$zj�)�K>pQ ��5�'��'ߠ��2*(���lY!zc�0
�'�\k�ǖ�pL:L����wt2MB	�'R�7�Ļ5iʠ �l��}8@��'��X�_9�T�ʡ�F�!���ǓQ� ���V�����(D'�p|Ȣ�3D�����  �'F>�БY�D¥p�N������?��O�`M ��4u&�̧O4���k���W�ID�4��B��0<�bH�Q���[1!-}҆K!7�[�"'@l a#e��0<���ʟ��	�����l��}Ҁ8@�؁���XѮ1�'T�����F�xu�����"��'H4�����(0tnРl=��B��L�m`���%�O˓3v�h�����y9��Z��]͆�7oMeM8�'�- N��A�{��I�2"Ȕ"C��X�b��{E�ɩ�4�b�����uH�%V`��K"�
j.����	��@&?��|27��� 氹�G5S��Sӈa�I񟔇�I&I��0��Q�V@*M�gc[� ���?�4�Ӭ L;�EFO�"�J��ڙ(����\�`⟜�S̟���q~b �1f�^`Ke�4Ac�c�&�(�yR��5I&���D�R<5��
��
��y�H��V.�bĨ�'> ��Υ�y���%|G^X�5,M� k ��S;�y2k�d૥߾����	���DIA���X���.X��@�T�}t�b�:]����O.�D�OP�O�'T����j*!tةĄ _=�/Oi<�q̌2s^��S��]F<ձ��Ԥ/Z:\���s_��R2��s�ƕ�5��	���w$ៈ�Iܟ\��Iyʟ1O�8�d�3hjq;�LH�&�*��.D���f�Ƙ0�b����%H�d|K$�'�Eڦ���OyBLz?�ɟ.�8�Ό�}���O�b�^Ě��'��'��<�B���)� h����n-��ðiO:��f�'JX�J��dт8#d�p�S�
�b�M��M�ax򠋄�?I�yrLV�7�|U`�!�9�� ��.�y�V9*8=0�#	,3� �H�����?�2�'PL1 b������h�N�MX���ҫl�����AC���j

G:Ÿ��[6R�u�������	0a��$ڣϒ/*0,lBE�¾l.�B�ITQVm)�D�w��ѐ&�~NC��-+�����(��[��s�+˿0K�C�I	\̀�'�.Y�XMH#$M�?��?��퓨)c�A� �Z�P���O�!!��ċqO��S�� ��z~�i�"�V�9b�A�]��L{����yBI�*.D�� #S��+�^�y"�� �k�ፇ6:���y��M	���D�%/��0�R��y2�Eyֲ��Ќ�25�p�%����L��(��)cL�*b�*E���"H`�3V�TsDK���\�)�3&.�p�_��PU�HݮB�Ɂ2�����e�*Y�@����O��C��sy�T棔(H���q�ːl.FC�IZީ1�f�,�[��ȯ(0C䉺I�
Ĩ��H? ̑�%J$!���O2lE~��M��~BaW�J��8B��Ũo8�TH����?)L>A�����I�SH ����g�4Ȏ�2��B�	� s�9�S��+29�������.�B�	5AF�XR&�4*�ب��P�R�B��eN�uR/�P���N�G(@��������� �5�ج��Ŏ�m��t��J"ړv���D�d 7$^ ���(ƨFf�	`��2�y��'�a~���|Hh!B��6$;����y��A|l9�e�c�N4�1i��yҮ���#B��.φ)cѡX��y"�R�hF�y �ޙ����w��+��O\�G�d��̾��`&��[2�M 7���?�7g�����'�����p$��
��3�S(=G�	��#D���ԡE��9�ER�\�]�`$D�p��I��R����WK	�}{S�6D�h����+>�8�C҃H(5��A��7D�d3 ��5)JD����m����@�<��)ʧ �Nq���]�^�qD�7UJ��'������'���|�����8e��h97\��4��BA��ybcN1n�Y��D&����܈�yr�O8
"�P Ɩ�A�E ��*�y�$Kd�8(rA�@�U޽+cNε�y2��h!u±�(
�Iq���W���Xá�����U���J�j�AR �?<2P���g�O*�OR�d �3}�+�����h7HךnО0�#���y�n�
�����n�hi��Ŋ�yB�]7i���)�m[�2�c��y"���bH�H�mL1{�����?���'>���R�I6(Ӏ�:�`W*e�8=i��DR0�?U��-˪�lD��QYP�ן\�	{���pD�	l����0*�:2���q`�(D�H��.��xh1�I̝e�v�&�3D��s�״X��9��H_8HKf2D�t��c�[���3�o�+�.�'�+�j��>�P@ȓL$L��G�B��h���O~�2��i>��	ݟ��'cH]��N]4Ռ���D
@ifU9	�'���l�5rg�=k��5��;�'C� �c��
7Q��ٰg�0�2��	�'B@1b+��C6��C�J��&!X�J
�'6H��J�.��)rr�N��T,�)O�Dz��mV�)��oӴFX��b�^)Q%� 2,�d�����$��>y1�*��X��N�MzS�!D�� L�
Uh�9w|1f�ƯU�8�e"O�Q
�#�sd���F��
Pk�"Opա� �t,�D���L�n��k�"O��3!L�:H�nt�@b�U6�S�|��,�U�t�="r��b�ւT͂|�$�˚S��9��l�ڟ���O�C#�G2:�T��%�,'Y��Qq"O� *��@ЀKD)KV��yB�P�=�����⅍ 6<�îK)�y��V�B�"e*UFԬ|teP�(C���?W�'�Q3�H	*rD���)+� i0��$�+?��u��T���0���+��9	�
�����K���r-��,�Y���u�Dq��6D������&U���/ �I�4D��I��-�"y�H\%T
 �Y��0D��@r�J�-�IYA�;q�9P�j0��U��>���D��N�Z0-A�Ќh)�O�)��i>��IڟX�'n��G�O��Iu� 41|���'���뗂�9gAJ�
pGX�!� �	�'�J5�d`�;g��!�G$I=^�jH��'Vؙ�����pBK�]�8
�'�@xbA�Ɯ{JT4�gd�WJ� �-O�Fz��)����y�m���<K5��	���	N��y��ԟ�&��>�����t�R���)�&,1Pb3D����:r�s����Q>��m-D�4A��2HvajC��%|(:e�(D��XGH�4\f�ɢ��:r<8aG$D���1�+��e�0�W/r�t�q!#�d�r�'��(C�'�25jca�dՔ�j1CۓY�Fea�����?a��L��҂��GF��`κ4�6�#D��H�η�X 1��ا� <�4D�P���{�d����/X��]`s 3D��1n�3ey�h2�!ƾAۼ!Yt?�O��	�:P����ǀ l cF�Fȣ=��O�k�O�ݐFL�nr����ؾ!(Y�'�"�'5j\z��AR򎁺�`Ȣe�'��ݱc̜�R|�w�:�`��j.$��B���P�AbЎҴV�tm�ȓ,'��۷i��p����$�˭EZb�D�� �'C���T�œZ�n��m�?���I7?��#<�'�?)���dч:��Z���&�Ԉ"��ܫ.!���d��Ư�_�v(�X�(!�
M¨�CLH<+3JA.Aq�!��	1E��@kE!3�x���,^.@R!򄔨g����`��<�3���l_��=�HOQ>9����2{��q�D���ȡJ'	�<�1n̆�?!���S�'SG~��$��:\�'�� ?�
���)������ʚxa��d%B2N�Ʉȓ ���`f��{��MQqoJ2\q�a��9/�qQ�*jN(����� ��ȓ4���+#h^6yR��Ka+�;���'����$B1��$�0l(e�H�e��D��<"�|��'���s��9��;ޠm��ǚ�]��@$"O~$��?c���b��ۮj�D��e"O���TcL��:�0d�Ue�����"Ot�� �N�����EG>�x�9��'��D+L��!p%/8R��z��z�ў�h1�,�iqn�`I�L������MX�<���?I�/��8��b���i��]	%���ȓ|'�Mk2΄���`��Q<Eh�ц�Ԙ���'j���x���%�L��ȓ#z<��Lט&.|؃�E�J���F'-�'<m��Ӆ;.y:�8�b�9o���	�N�"<ͧ�?A����ѓ�m3H�,x��Gnǉf!��<l���s���rWG�q�Xx���� �z�f�5 2Ր���,�(a�"O@c��`p�)&��#A�+`"O����퀰s�P\�"�)M��Q�[������ӻtU\9�	�r�V}�0S� ʓXG4lP��?�H>�}Z���mH)�7�C���%B2E�c�<��K��@:@A7f�(4�	B7k�E�<	��<F]� �,¨���Rj�Y�<���|��h1�fJ"XB�8�'��V�<9�R,[&�1�t�@qz��P�ɦ��O�����O���V�<~{F�tH�	P�jY3�'�'���>��;���ӡ��7\�'�u�<�I�>$��C�ω1l<y��)
t�<i@YK؈��= `ei%�q�<��(�9W��a���U�ґ�5�JH��x;�:eِ�1.��]ra�C!� MD{�n�&���nc�Ԇ�d%#%�)!�F(���O��D4�O\�
����;�*� S.�&tx�"O޵Jf�3|
�z'R&��E9"Ovy)�gą�.E���1d]�R"O���p�@�D3^��b ����5�	��h�zȄ�Ft����攐7�����'������4�V�D�O������i�+�\�N��l��a�ȓ"��j	R(�V.͑r��ȓY��1�(�";��u��6@�n��]zT9���d2��񦄵=����1�
��g��?ޢ�����'�6X�'� #=E��'[�p����Z�s�@(3u"��������O�Oq�,LS�꙽w�lZ��(4g���7"O^���h=X��a�)�"&/��S"OR����B�l<hd���\
U"O�9 ��P=�!y��ܵP��D�r"O�0�� �[����)�O�P�|�6�	����D�>�a��:d����ϒ�&:���^����@��O� 
��YN�"��Qa��M�H�	�"O�X�B�E�[-�rb  �ޥ@"O�d�e��\����͌t�&�!"O8ĪG�ĲoC���a2�@,���'�����a� H�3r^e�bᑦA�ў\F�8�u,:�H��Lp���F�,^~�(���?I�v�)˖��?H���	G<?�ȓAX�I��E 1̽xШ�N�r�ȓ_��rGݳ_�m�A�ػLp�B�I�P0��W�S׼�R*G(EjƢ?9�퓥R�<�5mєpf�`�j�l�~�D�%,���L��p~.F*�R=Ҥ����퉖����y�&��i߲���H�s�����y�BY�����\�m^P�ˠ �yr��/W���aFیi�ZIa�eP��y���>0��Ö:8;���.����$�p��(��y�AI�2��XKg�� �ΜHR�d�������IL�)��0R~`a�~�)s��ݼ)�B�ɂJ�2�Ks�֋�hU�@���C�I�l�yc%�L;=�2�+�B�$Pd�C�ɽCd04I�f@!T8�4�\�kbC�I"P�>9q8�U*�,�(�Z�O6�E~�k���~Z��d�*�5!UaO.O@�����?���L�(�a
�|�,I�vi��ǐ{�!�ĚS`��*J�t�t��IT*a!�DN�k���fㅃi��GH�[�!�N"�­p���$V�xS2Ǉ������O>����I�|�yq���'al��e�I>p��#~B����kjƙ�`��}'�"R΋�?���0?�6�-^KL����$�va�U��x�<yM�1qF����!c�h@#%a�p�<� &}��̓1b���te^-+��c"O����DybP��7�R/R ��ڳ���h�=H�C��S���B�J���'�
����4�$�d�O��P�8i�C���g���P�;(�����ƪ�:$�G�$7>�	e�7q ���Q��q���%U�����ƶy:�`��3��\ぢ�R*�q�f�1\�J���:�$<Y���*̦���-�5u�@��'T�#=E��JS.������6#V
�?���1P���O�Oq�lC���	1N4��TO�$
�a�R"O�u��*t�"%�a'I2q�n�f"ORl�C�M�2t��(PGZ9/؊M�"O�����S��<���3hd�hc"O��2�P )��bV�;�	�1�|2�)�
y���:��J7��+W�|��g��x�ҵ��m�ϟ4��OԀ+�X>|��l�a߄j�z��"O�zզ�>=� �K���!��Ċ�"OP��kԼec��4Du��iE"O�����͉�T���蒉�H�x�'�`�D\�,\f��SCćm�T����K>
�ў<��4�.��L)�ҍ_	d�@	G��>�i���?y�l�r�K n��u�T�����@��N����s�4��m�4�Iٮ$�ȓ+����X'`�a35m҄-m���~i���pgN�8�#��AQ��F��<ڧ��'%2��ڤ��z���0�#<ͧ�?y���d@�|��٠;D�i�W?6�!�䑺Rx�9�&�B�1�,+R�!�D�9qF(�\
2)[
�^S����'�x���L�DSX�rIцO���`	�'0��`S,Ǖ'T5�FGΔD��I�(O�aGz���M�9w��Z5���(��MC>f��6}��>���i}��>�u��$O�F�!Ǜ�H���0�B�?���?1��d�����(+���O�O۪��T�P�_�(E�iг/�J]i��d��h�����l���3��|*S� Bx�Y��dǙY8�-�6Ƒ|�'b����?���F��dʹI˜)0̾\�����D5�O���WN,����C�r\Y��'���A�@>_&Z���V�-�&D�'��ِ�'l��9O��6D@�0 �׵\|z�ȗ�O�,)n�$�����Eڕlq6��$��"~T�ʒ��y�+��i���	���<93.Q
P�4�%ɐ0Rz�:��i������OV�\�jlp��΁8��M����'X�)�)-?	�A:+�X��¢i�|*q�Jk�<��,D9�"lr�զ+<,�Q�c�'p�"�c�0)��<1G�;q�dCB#F9B�d�P���OKb�'��'Jp��-�-3%BU�umń#ߨR4"O��(R�<-��	59�ʧ"O�iC_gx5�#*íN	��ڷ"O8��a�
�����Q��"O���,Ű"$E�.� RH�P"�'7�#=E���"CE$䃲�U�38�X��T� �����W�2�'ɧ(��T���_+!����_��P3�"O�����mD�}e�������"O��g�I"'c�`�6+������"O���˘w1T��5iw
�$��"O�ͱ�(�Q�:�� 4Zd�U�P����DܿK�f����/S:d�ȠelA�A��X$���I����ɣe�C�(-P&��O���C�	�.����'�� .�#��B�ɻu����!,Wإ* J�>m��B�I�l��%z0�F,G'�՛���)O���Vy�v��D@�`��A�'H���'�h��4����� v�f��4�N������$-��#������e�)Zh\hW�(D��01h	L ������*6X�p�+D�� b� �D��J�����E���v"O�����,�����`F0�HK퉳��T���Q�V�t/�0{��}��Z��O|���OD��<��	�Fw�-�b��yk�e�\�B�ɨ
w�-�!DHP����V'ZX�dB�I#_T��'GS"7�	�3&��J�(B��1p�0�D��P�B-�fh�x9B䉂:6�x�7Eߌf1fe:�o҇L���dTx�����c��ڣL���3�hԡ4Ib���OP�1s�O��$3�哄J�J�X�f�B�`�C�I&W:H
0EL/`F,u�� �>?�C�I B!Xݚk�/#1L� � t�C䉨!i�CP��2�A$��N�RB��!e��x�B�J	3Gb���ƙ�,ʓUڑ�8�tD2}���r��3$&�:��Z�3���?Y��0<b�g��@��_�;Y�@b3ms�<�Q B�]jv��¤1�J�R��Hp�<y�f%o��Y��̗X��e\x�ȓ]����E�]�XR���لy�����	;��ހ(9�$!`N�#YE��ޙe��	���	~�)��R�@�ys�\���a�O;LO���禅&I"���Wg!+n�`v<��즡$���	V6���KW��<.-���B闇 ��I��~�ɗ���|�j��%#W�}�#p#X��E0�kY����FT���h��~�O����!�4mwJ �p�]-@l޹�W�g�do?���9Oh�1Q��h�vB�$,������J�JA�#P�%�Or�O;b��P��"�蠠Fs��3�R�ݦO�|�g��BҶ ��C������^�p�E�ɓZ9��'���'l@�zM�0�ٴx���v(?1d|�c$ ��'�А	J��k��锂[��Ucp�*���hL��X��-?P�O�s���??Y$�B�<��\�U�ǍqR�����Y^(��+O�}!@������l�ȥ��IB7jp�h
�<�H���9�~�KV���?�	�Ayb�	�]�(��d�ZiPy�0��mh�$�İ?��̸��꓌�>��;�#�[�<9��Jc��˔�n3�(��3B�IlD�����e18yq�b�nR2C�	�W��L�s'�]&Ҍ�P��7`C�	�>><��L/)����&ÓFaXC�	�y
(<�#擶8<��@�@�:C�I/��DI�T$����F.&
C�I"i2��O�w��d�τ��B�	F�,�@b��8_p$��ܳD��B�IZ�R�C�C�Q�PbP�h��B�I7,��r"��'����C��.q,B䉜L���QD�{�D�JP�՟0^"B�I�
82��U�W!Б�ňR�B�ɿQ1���-Dif����7�#<���\"}�*��]�̌��HǀBy�U2���:����F�2�TMs��L���0ɲ��*apX�����1=~�DY"I��0]�� ����� �C�/�\��1��0%Șt'͞�m�VY��-��3CL�{�ĉ:��0��l��S��6�@�+�5X޸�ʃlϳ*uj���,�����h�5 b|b�6(�����=7��)�r��"<�T� @��� �R)�`n�/s�����
P )萮��1*&H�p��1T��s�_�p$yb��!cdm��@�8�(Q1b	�u�̃CA�(gtly"K>��+�%-F a���g��P$�@H�<Aw`��N8��@�8.�>h�E��~�<iBL(�>��s ��`W∢Rd�w�<�㬀a�ƈ8���0Qz����r�<�T�׎.��2��ȁ^�,$b��p�<9�a�',�)��_��f-JVg�v�<�'��3PE��)qO��X��uz'OJv�<��	��d��R�X-%Ǻ����HH�<�b�Ǽ��%�ë�n�"��\�<��F�N��v%�uq�}���l�<)m��R|����"KX� :��j�<yb�P|�1c"��$H�jM��N�Q�<�@fS�mg��p���7i��-�M�<� ���C���xU�P�b@ {g�HU"O^���^->Uq�;guP�"O8Y�E"L�LhPoO_g�,k�"O8R�%��/r�R���~�4��"Ol`�J�5?�(C�됛 F�R�"Oh��L]�p�ք��1�i"O(��0I�jU%�U�ՑE�hH�"Oz��O��n8�ae�Xw�� 8t"O�1�j>)�d�h$�::�\�#v"O(�6OGN��1�)�4(Ph�"O&�Z�Ӡ3��1{ ���2T��"O ��` �	Ј:D�<(����"O�Rխ�9�p0�'�r��8w"O�XQդ��P�x��g�\=u� �"O�$b"�՗Z9\�� #׮��y*A"O6�٣c÷qK��Xu��+_uv)��"O�SQ��9��Հt�2"OX��L$BM��lhO|�c�"Oȕ�`��-��	 ���d`�1#a"O2��%�N#?��[�l��R��(2t"O ���o�9ql �{@��{� ���"Od���)���@�k���i�<|�4"O^�0$y�y j��~�`�"!�yr��`lŊ��A�����	��y���"\_��{a%�V�ٓ/��yB'��`n���a��R<i)��R��y�!|�b(�v��+u��2�@��ybbN�`:Ը�LW�g��Aķ�y�ˬ-h���=a��a��?�y�&ۜ-β�e`��O�: �׃��ybo�i�~ �4aؑK��)1�/��y�BJ�9⺼����B���%��8�y�1*��c�6�����-�y� �uU��m:֨����7�y���(�l t�4����)�#�yb ���,�J�.�0a�'b@?�y")��~��]�?���V����y�+��R�b���A�=A�Ԋ����yr��w����&�K�t.�+�y�oH�,��R钀v�"%����y��to~��%��gθ(CmN��y��N�5��9P����i�Eϝ�y��_)��-yŋ��J��Ò��y�A�4L�#�ܝ�� ��y�F|�u� ��t�T0R,ۊ�y'� ���)n�%r�9q톦�y2 �:6�up�/lc HBa&�$�y2)�.Vv@�F��-~�Z����y�B�(~�xCT��xy����#8�yB�=�"m�w�*_՜ȋa� �y2�Y�gO�\Y�j�Y�J�@H���ya�>{ؽ���'�A)0��y��7�j�q�kO�J?�`t�
��y�B���@ D��:20ś mM��y��!����f��+:`�I�gG�y�&��,�bE�w��05t�;�]��yR(U*�D�eO:u�1��#�y�k�3(������'J9:���y�E!ɪ�`U{���CO��y�!���̚��	t�|@��M��y"-ϻ"����b��X�>�顈���y�OW�^���P�o�:GR�Hi4F��yB���>�ʤ��,�4B�h��"��yB���� xF%6�B	�Ʀ���y
� ���v�Ę�B$�ԥ)�f�@�"OVi8 ��6pR�K�>2���i"O�I���F�,�l8�c�:|�p@R"O�8� i�.x��i�X�b�
�"O���2W���W�M�(@X�P"O6	z�
9\��ZP��$K:�}
�"O�m"��Ȼe���"�)d{�Ԃ�"OjWnڞ �#0�ҵudvHs�"O��A��֘;
ȡO�zD0Q��"O����!W�\;�MS!D2���"Op�l0"���1��O M�~ �"O� ��2H9���89�ԐSf"O��)b�W��0X�Bk�7,�
�s�"O|P3����������O�R���"Oru��*�zP�<�
�&tEJ5�"OPd1�N�w�J�ǋD���u"OP0�D6E��!Rċ!i�f"O<��'�ر{�Ђڰ
�mK5"O\L�B�J�sp��VK��t�hm"O�� ��!{z��SJ[�v1�	b3"O.��SJٰ䥸�nĂ(:�"O��ࣦ(H�V<x��V�xU"Oj 0��λkچ�ɦl�6;� 4�"O氉 �Al����4kN�S_�a"O�M�V�Ҟs��T��W8YAK "O$L�o҂x�6��〙I�1ڄ"O��ѕHh��0���ķh�N5��"O�U��a�"D����ˉ$_��P�"O�`�	ܴ=�ʳ�L#\��]�3"OT��F�+�)��l�*�"O��6+Kw���0�٬�x���"O>��q�.�p�+5��?�~ݛv"O`q�`W<<�l���>`�ZX:�"O`a(��=y����D#&����"O8|�ׯ� I���ڠ�V�?���8�"O�T�P_��"���0k���v"O����[L���1f��a�"O����+��M��895�y6Ʃ`�"O�J4h��n��AP�c�`'�Q"O�q
��֯Rv�|�g���"O���� ۳v�,,{�Y�R�8�"O�Ö�����8T$*����"O�\�d��L��l1�d�>Vh�]k7"O��@K�<k��a$D�-EVD��"Oؠ; �?��,Ţ��+D�j "O���F��X}4�H��<v%��c0"OLl�ueS9F���RkA�D0�;�"O��aF���LU�L���<^��p"O��0��W�?$4���+Ѣ=�BP��"O�D�s/9$Z���%��q�ݛ0"O2H[�b? �j�;�&�Lmh#�"O��"g�Lˆ #�CO.\N�;F"O��)�d�*J�tAT�ZgF���"OJ�I��C�6�Pxه��}8
��g"OTZP��)h&��o̱)�4ằ"OuX��/Ww��(� ��>�P�Ib"Ox����,.pP`�� Ա"O�-�G��+��"��[�ԕhW"O�\�����~�8=J�J�(0�Tѣ"O��K%��z�zD���N(���"O�L�p�)!0VA�Dh��-4"Ox=�Q�N����RG?ZK�Ч"O�qhVI\�R*J�buE��$Ap�ڡ"O(A�`������S��`�`"O� �Y{&aO�F��(��ԩF���A'"O`��TD�1qfxY{'��Z�1�%"O�T�e9J�vi�g5<��=��"O��"A���S`d�bd`�XWB�#%"O`Q�N�I+���hF�1��峓"O�Xx�+��q�@<��GZ�J�,�"O����-�J�65��� "|x4(�"O�< M	;9�̙��Q j:0�2"O��p ��\�����)/��@�"OFij��� %|!���X"�Db"O� ��J�^)JP�e��+�h@%"O>�4�SP�ᚷ���I�p%S�"O�q�WDQ9K�p�DeQ29 ���R"O �jDB�-ɳ���7����f"O��+�2�0	��V$	��0��"Ox|ZҤ�R��"�a�#�l�۰"O~�Ј��@Hk���7�D���"Oȵ��܇o� q��/�_���I�"O&��D���!�|AC�8��u�"O��p�ѫ.~��2�N�%{v�;�"O:�3 �)!𨫲��0z]�"Ot5SHF'jޠA�D�l�ж"O0 g�m�n�0T"�8r��ur"O�Q����V�Y�$k�:a�tL�"O�iS�ڈ&� hr2�H�V�B��p"Of$�LP�"�v}dL�
{���"O�&n��e��(�G�Y�	µ"O�D����;|Nq��&��Sq"OҘВB��/��u��F�<|y�"O`��s���/·>��7"O4D���5J�x�0�`��_���v"O�c��� ��S m�}�@Q��"O�����QHhJ�#�e�.�� c"Ob�CeA�!�2��F��F�: ��"O&�)�"�r\0�[�d���Щ�"O�p�3��?<d,��D
!F��x�"O��N�,��lp��R%s!�\p�"Of�:Q ˙;-Z�7�_%�cb"O:܂S�ɷ]�w ^�$D�X!"O�,�C	��>�� �IL��P��"OD���L�Q&��0F� S$"O��ӄF(&�uȦ�����z`"O��q�'fU�#����� �"O~��g�\���ӂ7��;�"O4��¹��)r�! }h��G"O�I���G�r���h^��"O��)H��5c7/�S&�A��"OV���A!*\��6�MzyP��p"O�E�s�Ϊ3͜�*��ݕsr�y��"O������0$���R�=({.�P"O�`�q�֝u�Y�2G��Dz�(�"O�����u��"aM�w��}��"O|���m+1���)uZ��ei"O<D��aϋ�a���G�Xq�G"O���k�N22ǈ��+�"Ot��3ʐ2&�䐣���"`����t"O6�xѭ�0K�.IS�/E�)�hp"����zt��͛N5YvM�^i�'�����[l��E�B�N)�'��g�*ZV^���\&|�X`8�'�ܝ�ơ/t
=�c�߮!����'��`�3�e@L��"n�i�X�'B���t��=W���#aoG�
G��	�'��M!�"ПLN��0�>L`����'�����	o_�{�.ԏE���p	��� �T�4搥!��Q��='z!�P"OR������kH����>3|f�pR"O�]���S�.�>���"Άdl w"OBx+���U��dK�2PT#"O`)B���UM<u��ȓ�1J��ɕ"O `�/��y`����|��"OL�������bv
�m�dt �"O�M�A���"�pJ�&	���"O��SEFN'�Ը��c�a�:�P�"O(�2e/՝
�,�r�kP��b$"O�4�S"Ӂgd�ٙ���unt�"O�u���E=Y��o1p�-�"OjPX�h�-\��]��i�@O -�'"O~���*E�W�di��/X�6D�a1&"O��h5�ؐ?�zՎ��\�r�� "Oq0���"p<� �������Id"O��+0,��i.��Z"E ���@R0"O,����!7�\<��AB�u���""O��(�KÙ[�fQ�R.\33���"O~�z4�?S���c�+�$lj8�U"OV1�à��x\!%�#1��A�"O6��_&s#B�u��6�"OZUJ�`J��tAk�F@�Mp]��'sj,��b�,Xb�yjg,ߖt^�Y��'��X�����Z���
�LB�~;r� �'���a�lҨSq^��q$ÈHiLPa�'�)Z�hP����4���.!@��'�����њhQP�2����'�t�)D�Hj�%�s��7*c.l)�'.TtS!̢ɺ J%
\q�'A��s��A%B�ATj�.��a:�'̩C��t���┫�� ]�,�	�'`��ǂæ5�����W�.P4�I�'��Lծ�;�9!I�)[(@�'���!���FgB�|�j�'f��+/̥VjX3�#�9�P���'�<��C�_�x���gĴB�L�'�8�@T/:�D���.�K�Py�'4Π# BѠ��Q�C��-0=��'&��1����oI�%�Ȑv]��'za�	�ZfB�����|��'���B�"DL�9ϗ�M.$;�'w���Ứy��С挒q��r�'�ZMyƃ�O���a`XY��T�
�'
�	�q�Q6�bq@�Z�[:���'A�e���<����3���pX��'���F�D����2(�*=-h��'����" R'N���B�7�l��'���CM�8���+A*�%
�'5��AC �/\uh�#Wo����'G���N�>jװ�4��k���S�'�\� �ZC��-�h����'�b]ص��z��k��ϓc�f��'��)!�dG25�=R���4\Z�'����RH�4l'($A��S�"��:�'�`�A�'ϻ}(��4!��LBI1	�'i�*�W.;�:%#�G
.H�r��'��a���	!d�Pr Ʉ�ډ��'��u��&�)a���ʆC�kf���'l���G	[�=���ڑk�2�n(��'N:�y�	"���B%s'&�k�'��	�2م	�P��p�^��X
�'&pyO� �"]�!��H�����'T~<�Ύ�/{"-t�U{��(���� tlu�L3q{b�#Q�@b�2"O���Ưv}4YB�k��
M�)�"O�� ��	4�>�EhM�y@�m[�'XV4XtE�2c�;�EC�_�fIy�'�� �鍲K+\�@�]�
<��'*I#�T���V(2M�2)�
�'Z�b �?�8f�V�Kj\j
�'�:mH&�M�xy���߼RP�u��'B���W��j1lLm�E�'QșQ皈R�vY 1d��.��ap�'~&i��,��ԑSuF��-��J�'���!]);��Q�']

�	�'}Ԑ�����@�`�aԋP�a����'ȡ��N��%�GmZ'`����'yؼk@H
�1�`-Br��8�{	�'E�ٸ���"�M[%��.ZJ��	�'�"`�Q�[	j+�� ���"AH�!�	�'� �HB�)<y�@�W�7A�Dlj
�'�jq�kY9$�(���̗v�$�' l�rO�&-|����A�;h��s�'�Aȷ��7utB�!!�ܞ,�$�@�'���C��^�~�H�bJ�$SF���'���i��_Z��� ��*/�v]+�'~����A6� h{ B�p��)��'ڪ��]6�"�X�ϋ3@��'��[P�T�s�	sǊ]�4t{�'2H1s��A��qҫ�*Sg��	�'Iܩ��_N�xy�'@HE���
�'ۜ�;d�y�\49 B�0}��
�'�9� f[i��M0e_;dxP,3	�'2����	F�8��B,U��|	�'42 ��TÚ�SE�Ɣ
d� �'w�P'%Ƀs��|�g��9�eB�'�
��
�I3@<�I-��a��'��Œ�JQ��`C�1[�L�[�'�xa�5��t�D���^?%G��y
�'��b5K\�5������#l�$��'{��9��'�z�+ �Ȅ:5�e9�'�����h	I!~9p#$�03�%��'��\�����}۲ˇC�_���'�܍��h�{場�WLėPǶq��'#:l��u*oޫ2�XE�	�'T����o׌$��'R�*���X	�'ǆ�Y�KȳXdlU(�`ɺ%�����'���0&b<h��ㄜ�"�ݛ�'x������?d�R��e�H�@���']��bǁ��E���Zb�����	�'��2���z�0�T�P�W�Ż	�'HT�A���*WH�t��R�I�~���' ̬���K1LĞIITf��}M4���'s<�rk��a��Y�ǥ�@�4A�'�@P�N_+F��F�7A����'|XA�\%9�|�Q�ͳu{z���'5<H"�	C�!I2� oSԬ8�'�H��擆-8ƴ{�΀�l��%��'������م���nD�`�~�:�'�u��'�E��mRR���l�'Ih,�Rj��S�)��D9}G��'k�īSl�(b:�)���:�8)��'��4��Ԁ#8�1�b��N��1�'��K�84 �E`�$ۮN����"Ol�q�čGv0��ʆ� � Qc$"Of�!H���	p�䅟Y�
�!0"Or}�7!�Hg�c���2��}A�"O� b�[P�
8x���ʡ!�+X�^� &"O�%�!���xl�S+˶D3��5"O��$�3f�䪰��Q$:�p�"On-b�L�"�*P����q6H\P�"O���e!��az@�Ŏ/"�H�F"O��Q�E�8���2��ز9��"O���F� /%C����ސO��zf"O2�J�.@��J�1�Q�l�B�"O4� ǋ3Y׺����Q#t���"O���Qʎ�(��� '��~~�8D"O��:3 X�%˸��P₄u4���"O�pR�Ɠ(p�����>6i���"O(��`��&a�J�St�Ҙ#�Nxx$"O��b�G�	Y��Y#I
4�V�Q"OFi��/$m�#Q�&�B�z�"O8�80i5G������Z���"OJ���'Y�5vRp�2��;w�x��"O�e�w��s4ʩh���7j`�y�"Odh���O�XheC%��f�Rq"O���N�V��ʂ"C�J8�8�"O��0J¦H���T) ��(;c"Od����[?&��Dt�-,�����"O��YSG�3�@ڕ��!8Q^�r�"OR\�"j�!Ǻ	F�Y�p�pm�d"Ol�CF��>�ĉ�a��4^nB2"OV�@��A=Uq�iu'K)x��d"O^�h�2��hs�fL4_A���"O���4�V�Sp�T�EE�pm��"O޵�W�H�>���ۀA�]���"O�`XfG�=�
�Co_�Y��(1�"O~��U��6_  �,��~V�"O��s!��'��<Yc�M�Q �"O؈(M�=��Pea�<+�!��"ObH@u��$V�xѩ��&uDp��"OT�B��	N�|��N�O~�	�"O��外�S�֙6�SPK�Ѓ"O4�x��;y�&�B�d��5���"Or
��"^�H,��E�.~��`�"O~�5��6d�Ѐ��[�ʥk"O�d�Qa��S��yP��'���Q�"O(��Ė!!!Rͻ�A�s�:�r@"O�p�@J�l�*Y��/�
����"O�q�����A��&&��e��"O��7M�,�p���E�p�D0��"O,�%&
�4�Xd� �U�.�&�j1"O�E�Ŭ��S��� G_E�~�YR"O��Q.�%�n�8"�Q�o�Ƽ��"O� �eڇr�~���� =��C�"O����ޫ'����"O:v:&�Q�"O���UH��WB��tD�)H$�4�"O��H�W�@��K�/D�=p5"O�����L 2aI
��<�|m��"O��y@��s��!`�(e���3�"O>(2H�)��L��B4O�Ҭh�"OҌ���B�PI9!,=Hoef"O�0W䛀H�F�Pp@�ZZ���3"O�m;���+[�B�s�kU�T����"O"�� ��ԘZ�*��L�ٗ"OtɁ�mM�rM(%* ol,Ȉ�"O �������@Fׯ	���;%"Ox(�0���"�4];@���;��������o�l���G�!�4x���"��'�LmS�դ�05BA+I��ح�
�'�j����W�Z���BG����'��x)�"��;'P�1���?'�h��� �jŹlΰ��!�I;@W��v"O�m�d̙!<NAp��:Fv)��"ONp��.�!7���9E!ج�0�e"Opp����r���4��s"��P�"O����i��\!���TH�+r�]k�"O��	B�*ph!G�}�u�"O⩛���w��8��]	�ĸ"O��[�BX��Ph�$�m�0��3"Ot�V�C�(P]�Bc�c���1r"O�����[���Q"��dxڈ"d"O�$sыIg��`��=
d��B�"O\Q$��2D� i ��.pZ�R�"O^U�"K�u��P�� BX�`"OZ��wR�6�Ƀ'#B&AZf"O^�ك�b�b@�#!
�'+0��"Oʌ�b��8�$��> ���"O�]�@�#/(P0�:8�0Q�R"O������*��|���X�9:�"O���/�� �V�1C"O4�)��n�[�`EmS��xQ"O�:� ��j�<<���#�嚅"O%Ň�89EM\�r���@�"Oq�bZ./[�HA��R�XA��"O��yH'W�|2F�^,�Yڶ"O$A��/3��4�7㑦j��""O�Ջ�N,l��G��u0i�U"O��҂�6NX�gAC-M$<�!"O�u+#Q8$��p�Q*ZN���"O��)��ň�!�GW �iS"O&�jvf�'EXx��L�s$T5��"O�X�!��е����;x)�A3�"O@���'hE�t:��7J#�IH�"Ot���N�IQD��$��m
�$�1"O*t�5�	7|z�Ű�����$"O|���D͍B�b0�ւZ,<�M�q"O&ũ�؇m�|�$@�Ht��"O����cx#P!H��� t%{q"O�P�է�)V1�C"0����"O
�!�O:A5N�L��A ��d�<�ERZo��e��)@(<�`�b�<����2ѦA�gȁ;N/�d�E�F^�<����-Y0�����EH�öM`�<Iw�Yw� �
1��Z����d�[�<ّ�Z�j���&0�b7i~�<ID6
����DEɤ
��q㦝z�<yE;/�T�i�$��}Ԩ�I�E�]�<q%kL&Jcց�Y�L����[D�<�"
�4"X�Yb�Oӄ����c�u�<��=tļZe��>p�I�[X�<A̫Yx�5���/k�M��*V�<�O�0"��]�&��eHAi7!�T�<���� 4�ݠE̡N��5��F�<�ShE�n_�
%�6
|�{d�k�<qюD��D����\�F�:�'�d�<1 ����9�X4�bС���k�'Q?
�)I(=�`ЪL�
aPz���=D����Ȳ�|9�4
�6+�9�$�;D�PK��<�"|s¤ƴ$�x�@d�?D�@r�gP�qUr4$�`������;D�	�f��`�)�(J���15F;D�h h�W>p�+S+O���y4�:D���)��
m�&�ÀYU�|��h;D�̘�oC>��ӕ�^���h��&D��y�.L�w��S,-��1Ҭ&D�� @�CGΒ>���T�G-i��"O$͂���z5���H9�"O�9��U1GS<|��`�7i��q�"O� ���Ha��K֏��}	�4k%"O����:3�H����"����p"O��"R>C���x#�!Dʎ���"O� A4iɱ��=�u#�f���H�"OLt���M"dy�A��hP!�h%!�"Ob`�w�@&�$ �5��5Z8����"O��c�/�.�bH;�/�!S�`bP"O�q*��,q�`Ccn�LCPI�"OQ�U'�,#��(�!��G��v"OT��TdŲM���r0��B��[�"O$)�3���q��,y�@��pC��u"O��`�#|b��/��N�Xp"OT�j&/G)5��a$NT�$h�j�"OD�� nȥYT���r�Y�k!�t�"ONe�+�#)<�1� .<�8��"O֨���Jш�����T怢4"Ov���$މ?���[�$O�,m��"O���t�fj�4�a�J8�hd"�"O�K�^�o
�ͫ��HUu���"O:�b$�ƥXC	ԅ s|�+�"O�	���Ul�)��G�MpL0�"O���B�2�b%���Ū]T�ّ"O��Ê�h��zeʑ�qW�Ū'"O��+'�F�t?�p��k��I�Z�;f"O�`����f�(�k�'ОZ7����"O~$H�-ÒFN��fD2Y;t��"O�*bgZ�#eb�S���s�:��"O0equ	Ku��(��P�,�� �"O"�����(�Eт	[��"O� '/\���90tA[9$yʔ�V"O�3��%[�� C@�g`���"OE���C-h�183*;_�1��"O�Lj�n�:��x�5�e?�U�""O��Ȳ�K�yL�
I��5ȸy�"O�)x'Fɛ`R\�h���V5����"O�X�1�N�\���B��G>�	�B"O� �r!ؤ���nt�"O��Q��F��y��

VP�!�"O��YbO]�|,��;�G�]8��Zp"O��pB/rC*c@�j�||��"O�YeIY0C��lx����$<�c�"O��0��KU��U��)1�\+"OmY�^᠔��хh��1�"O�.-�>��ӯ�OP:u"����Py"�ց-�j����
E�b�Q��KZ�<I�-s}�}�D�]��p���V�<�6CQ�;l�У��+~6�0�jYi�<i�g]�K{F�X���[��-Z�<� L= �lQcs#��:���ѵlXQ�<�0(#b8�X��aX $ìzr�_T�<�A,�K���Ҡ]�) �Y6j�P�<��F��Px�y!M�Y`��N�M�<Y�͆M��$��U���+��1D���s�F��ˢ�Ӭj�ȘR�a5D��� ުw� 񂄍Тi���kw�6D�:�g�vhLŘe���fc� ��9D���Ɔ��~�C�'s�Uː���yr�%�:T�T �&S,B�@�W�yr���V]ա3�,_� )�Ŏ�y�U1�6��f�*{����G�7�y�*�dxi��9ykv���M �y
� �}�r�32L~)�+��+9֩s�"O�X�eaC�*S������-J.t�!W"O8iXt]�R�2�R�)�����ac"O�0��DP����"o_L���"O�Q�F�/J�f)S'�4Lvh�if"O�y���D��|���T#qj�أ"Oh� &��jU�:A�� Ag�x��"O���E��}�# �2G�*�B�"O�+V�$ ����3��d�`"O���I|"p�5M$1�*d(T"OV���� )��1��)�*��"O�I ����.�2 +S�V��Yx4"O.|S!�E+b���1ʋq�t�*5"O6�k�ُ,�F@�R/D�&����"O|ԙSlO�oB9aڅ8�ZP)�"O�JTIU�@�����`F�p-�y�3"O����ھ�\���aC�(/0��&"Olժ�ӾQ���2��],��H�"Opd��@�l�%)� ��!:��"O�j��@g�`�ѧ���QPz�#�"O�E7��Ba�	!�Ղ����hL!�ğ&?צ�w�Tz��	d�S�`�!�Ro�^���A�=d�p9SaO?.I!�$֑"���A�Y2)ZU���Q$?!�D@=l�d��R.. ���cD�!X�!�մ�H����W�f�r�ā=S�!�Da4YٵBW�C�2���d
<�!�Ĕ��0�-��0����}!�ߦ ��� gɑ!��XD��2!�!��+-�����=$o�D�t&�:�!�$�t�j���&K>cM�!���@��!�:pk���SK��H��#��<!X!��RA�$��S�PM�T����-y%!�D�C/
�@	�-!�H��/!�d��B�pZ"JՕ:�k��(j!�Ĉw �����\�|@��P?$!�;}Rp	��>8-��SEN�T�!�ď<^��1�ȟR*v�y�C��%[!�d� b;��B��8.1b��O�!��1H8)�b ��rWk�59!�ڴv/\]qE�F�!ZR�qEH[�I1!򤂟g�A��L> A�Hz2g��3<!��>�Z�����<=0�ك��}4!�$-2l��Fk�$,��	��'!�[$�\�p#״<�xB�Е)!��g���آhƞ7�4ٱ�D
!�$�4Xޠ�Z�M�j޸��"ə'�!��C�3�Tx���+���v`�	,u!�$VXQp ��ER�I~�R� �]!�'Dz�9�C͕ NK�.�>o�!��	X�y�T���$l�7-�6.�!�dK�V�^ࡢ�O t�~��W��1c���Q2%����G*� 	�y�ƍ�K�\h!��Q��`)��y2ɐ�a[4aR6J��F�vQ�����y�$]�vu��1Oq��j�5�y�E��9���c΀�Ha��⓭̲�y��~�4-�K;O��T��y�X�dfDyh��+�R�+$��y�)X�T���H� �+�
�yRaTv���n�a����oܱ�yRV4�2�Z7	�V��%*�yB.ѝC*�;��ǊK�hA D@I8�y�Ő�..��
)q������\��y
� ��3�ˁ',�|��T�6��3R"O:�20���)��H�#��/�
�"O�;��>.0,Д
�D`r�QP"O$	)��,0r��
l��(G"O��Rq�Yte�e��!Zv��Zs"Ov����F>Ґ� ��Y���1"OB�Y��M�?�2�;B(G;|�ȥˑ"Ot���n�Y�T[���L���5"O�١�� �*�U&"+�vh!#"O���fQ!�%Ҏ:��ܺ�"O �z���;X\^U
c�T�d����"O��zq�!��U���M!p�*y#�"O^�[�� vv ��l�b "O"��VKC�_�Dp�2�K�Y�}:�"O���G!CF*``&lN�&6�� "O<��mBi���딵 ���v"O44)C�w��9s�0���C"ON�AP-A0{^�8�S��xMA�"O(1a %��l�Y`-���D$b"O�p�%o:��Qe̝�n�%qd"O��� �6y&\Y�1��#��4"ORA+�!9�୍�Kj���"O��R�&O0מ`�u��!Q�F�@�"O�q�b��dx�PBʨ)��Ht"O��k�	E�8�<�B���9wԆY�"Ob\R��Pl� 5%��^)�"O����":,xH����5f���"Oz��f�Z�~���&��j�b2"O�P�"��t���@��U�I���"O�	�ĆWdI[Ч�	`1tX�"O:5���J64���E-|�
�"Oj`Ñ�ٛO�~m��E8���	�"O2��Ȕ)��i;�jJ�{��2�"O���"CB	"�U���_M�¸ s"O2 
���TM��p�_<)�H�&"O��A��wla����>�@dc�"O��¤,J9{�Ta /N�mn�e"O�E;V��R�,-ђ��eHL�ڣ"O��b���AK���N˨6.�a"O �z���i�t�W-�}��l�	�'0��j 
'"I�0��k�D�V1 	�'PR1O<I.�۷�������'��؋ÃC�y���C����$��'by[��� ��y"���8�2�'H~}�r�>z�����'V!x��'fl��}/����J�G��p�'�Z��dF�c����!K�;�L��'�ƹ���ڟ?}H�"�9Lp��Clli22E�#�Y�����*(�9�ȓ<@H���;#<����@=k~�U�ȓ<z`ј4@"���4�Q5Bb��ȓ4�������7~�&�ᆢM*?��هȓ	�Z)���$H�Ѫ�z�4��q:�-��aH�h"��b���-Ņ�K��1��N�F�{����p��qɦ��Ug�?`�]v.р��Ԇ�Lr��q%O��IZ��G&ZO�цȓO�F+�/E��¢%D� ���ȓ~Z
(%`�:ak(!��#[SX⑆�5�`qp�++ʹ��j�	�:��~v<�"���j�t��!C�X���ȓL�鲖-�-d� �va������'�.��6S�5
Mi�^�`����ȓ1b�EJ�'JX����P�|��S�? �I�q��0XX�QE5lL���"OX+��ւ0�Q�BʱpiL�""O��e�O�8�|��N�{��A�"O�	�p%�
�b@��o��`-.� �"O4aZ��A0L���mF-_ ={"O�H���5��"��%��uh�"O��Q![�b�ܰ�UJY)b|�9�W"O���&����p0�IY(5mX�"O�=��+��TX萦�Vtcj��"O:1�f�-��Y(�'a��z�"O�,�aN/r�H!��ՙb�B �"O�lpvjE� `��pq́�|<:l��"Op���ِ[7��i��4e��q"O8���L�7Ϙ���mJ(<�^�ҥ"Of�y� �4��,hcmW�<���"O�����U�^$b��ј /nt�1"O ����T@�PY�F֛m�<��"O4��)��>U3��C����iD"O�%{훏=J�����d�s"O��@��(OB!�G&ȚH�B�"O�Y۴�A���t'Q�~�Ȓ�"OB�i�nR5v�"da�*/��諒"OZD�%X���@��d�p���"O�ȸrm��9?� ����3"|l��G"O�ȉ�ňu��Ԭ�1�"Oj0�A��0oS�A��A|�4*�"O�����)�
#FL�.�.�S"O�d���?�jq��Ŋ�M��tK�"O��	#N�o��a&5yb�R�"O<��/�jlag>)x�Y�"O��gm�t�0&\�J�F��"O��J4��X�"4�$��t��!#�"O,̻Q	;TRL$G>`ؼ��D"O�m�U�ԓ��5
�Ě�?r.�!"O���6��lԮ�+�$?��"OB}���Q�mm.|q6F�C��9A"O|��d��{٘�C��R�R�Z%B�"O�d۴A^�K�q"G� �r|�"Om��6���"������8�"O�%�G�9"�^��W-��N���B�"O�р��O��0�T�T��"O~l#����$�j� �P gςD��"OT�0�(E�r%z�Ȱ,�/Q��{�"O>����PT�ʤ��"F|��"O8d"�bJ�h�*�V$R#�$
"O���0�. �4�#d%�38����r"O�<��A;���:"̙`��Y"OBȑ0`�7/����d���)�"OB�C#N�^���֧S�4Ő�"Oh���
�ۊ(0��w���"O~�Q"$4~TY�Q�]�� :�"O�l����?L�ģfM�f�~��"O�Y�L�=5'h|0�,ճ4VH�T"Oj,)��_�@�h!�U��7>���"O���@}:�P��R4��9�"O�}Q�\3-��}C���S�E�$"Ol�H�VFLp��Κ+
�#"OZ1j�%��qXX�0ЏN�l� �"O�x ��I�"ۆOL܈�5"O( ��	ӷ!���� �O*��Q��"O&�pW�H�w�C��k��RC"O�$�V	^��,�q'X7Β�9�"OT��`����Ԓ����x�6E"O�p��i�hÀl�$��$/@P$s"O� (K�äy	�%��W�`:l�I�"O2�SԮɉ*�X�X@`�.9�<�"O�T�B�B^���1勨[*�IpT"O,ȥ�@�JZYB�uh 1R"O�EiTH�3c4��aaB#M�%�`"O��;��/C��,��j�08J�`1U"O�tJ�흠|�j��Ɇ=�Qʰ"O�YCgȤl�|	P�MRB��@�"O<�@U�����O�T��U"ONTD(��f�`pB��P�I��*b"OA��*�O
1�+I	�D"�"Oz��p�Ӧx�R8���T*\���"O��O��1����Ôx:��"O����-Oz�`�fb�!9v4c�"OȄ;&/�h�F��"쁍{ �y�"O�+�ȉY�\`rT�3\X���"O��'��?	�!1aBP�0��<:&"O������a���BG�[��I�"O6)s׀/<@��b��|�~@��"O~�4o�<��"@�o����"O�L��W�q&�\..��%��"O
�+��ո/g$K,��V���"O�у��
�P�ؐ3���NuH%"O~��0#�0�(l@��Z@p�,��"OrL�N�Ao 0��g͊D��R"O`�	F�&(� t�D;��@b�"O|EIR�O!/�(Q�p�Ȩ�y�F"O�U�&%O� ՌE�'C!�=1�"OH�2U�]�u�2�	�Ş��D��"O����X�4�l���$�& �"O�	�2i@�Vqf����6�@ih�"O`L�v@�8����*\@�S�"O�!f�I�"tKߩ\�� 4"Onl�ˎ�^��j�'Bd1�"O�=��K]`ae�1(-��"O�D����+)����cĦi�P�rD"O.!	���`��Qb0 ن����"O@�1��&!XeB�� ��Aq�"OV49�;��Q� Ba�}�f"OP-)�L��N�F�E��AD����"Oޅ	��D�o�T̹�f�@����"O���A�4c��hj���?n�X�"O�)c��:A�x[��M�W$l�"O�e�X��L��#2*m`�"Oh�Bq��1iKʰ`R�#qU��"T"OX��L�j�ʔ�t�\�PT��S5"O����+U?�vd�T���c��J�"O�4��?W��2�mݮy7��j "O�)A$�&),.hra�G&�(M��"OFTZ��(NSx�a�����JQ"Oڥ��j
z�|���E�U����Q"O�P�(~�[�V�m�:I�"O��%���
` �A�kd�1��"OfajĤB�~��Q������[g"O�p�b��b��X'h�c�.��f"O�16�W(3q���a�n%\9b�"O:\A�.ɹkPޑ��A &,r"}bd"O�Th0&�V�h� �'1`z��"O�� �� ��pBs��W��U�6"O�-����=F��n��fʸ�$"O�$�歋/R��ؓC�~��B"O�`g�&��y!��/8n���"O>��R��+���X#�VY|��"O2���"�7��)�6��65l%1�"O� ��"���1��a`#�5Mvd��"O��и����p�A.%����"Ob�a�d�R�պeL�*�5�0"O�`�Qlˠ&��ps�X�����"OrTk$���=����f��[�D2��۟��&Ҭ_s����r,�Űw�W�nQ��S�!��?�]�P2H>����I�6@��iS�U$#���XE�=���Q��(h.d �!잙V�8�QFS��II�7@�{S/Q��*\c���e�'M*iI���?I�����i�����紴{��	R\�����O��Op�d9������m�yI�!SgFiu�d�C;�O��m�ԟ�n� Z�hd$D=�y�jM6xۼ �V�i��tbc��ĸ<y,����Ob7-
"s�h�OO="���&�(\�丰a:E�ph��OD�'��<�aDׂ3�`D�"K {�"(H��Ϧ�������IT7Llq���3�H�kl��x���:�\`�E/ :ݛ6/��?a�����'�?7�@8{�H�E 1V�Tٱ�â@����O���(�S��(T�J��~B�\Y�$X)Z�<Y�id�6m)�SϺ+��:oM
1j ��84����L��I�s2��ڴ�?����?IO>��o���`�)��k�,����Qc�����۠�5#�O�1PUke=p+MD=x<�@v}��O�o����2��xb�7'Q����"�ype�`�Ԁg6��>/D���OXx���	���'�����ڗ�~!'щ]��y�5n*$� 0ףԠ|8�`�Y/#��� oӄ7-�Ǧ]�<��?ݕ'�,-sr�F),k�iæ�u⎍c��U�����'m"�'ɧ�4�'zE�.O@��)��n׌�*��dc� ���'�� �ir\��;��C�~���I����t�ju���p�����.\��i��(0��P�z��E�S�>�⑁�N��@��h�S���գ,�>�����%bۄB^��~�A%�S�O|�An�W��y���N35���(�'�x6_צ�'�J�K�f����.�)� w�h�3z���We�33���?��o5ԙ���ʊ6Z�I��x�O����D��w^�Ԛ� ͟�JT����H�N�d`Z�.Գ*yj��U��ŀ �J���Ϋhj@���HO�����'A��u�B�$�~�AA&<�����/	4�Dए5n"�4�|"=��MI�(���/p�<,���s8��Xش.���i;��A�[�����敺z���'���ĩ>q(O���<����e� `�4+������T��z�iT�Q�"�x��'��	>Tv9�!&Xk�61�@$P=�7�F�PW0��Q�U>?x�)��̄�H-.��%��r���¤�}Ӏ�P!�'�op�2�$=���2WWM�tE��'�
j�V��T������Oy�'��	�M��4�f)�7�X�Wh�����{Ӝ�,���6M��"��+���7���׊�N��&�ȅ퉂w�� p   �   �  �  �    B$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�U曞@�VM�P������@��P_`���'4r�'d�|J?��f�s^hy�&A�x������ b�8�`XTv�|2���,�
�*��ڹz7"a��iRȖ:[�Fi��	�[ڀ3�F�\l����S�
��0ɂ��O��d�O:�d�<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&��|�����$��::�i�V�%C���e�Ԋ!�lK��O4�$�O��d9��~r"&F�L����� �45`� ��A%h�d��o�&=���1���Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�Y�P�{ � T�>�@� D�(1! " ��Eɵk��<�s�j �M{��$�~��A�(���4 ��7�*��2��y>���=���O>˓ I��"��ߣo��u�)9?Ԡ��F��r����y � ыU6��ȓ~�p�k%��^��1� �
$F��ȓN�� ��啦 jN=H�Aއl�І������(����� #zy�q��K!�2�"MF�����X���KV�w<�%2�M_�I��$�OD���B<�����J��`9���)�!���r�¹�P�D*/���2!�ah!���#S_l$�f��dQ�ݒ��߂*L!��F
�L w	�zE���'�@�H�x��#���P�P��Sap��M:L-���J`eEx�O`��'=�)� (仃'یBx��"���6�˰"O�q@�	��@�aKb�1h�Lm�"OaP����`��\���3��"O���lr��-�3|�z)�u"O��vJS�-��H+A��usp	A��>i��)��1j�L�B��ΥjՈ��1��+���'*T��d�'7B�|J~�A��99�p��G�fp�3�C
Q�<Y@��d�f�B;R�&D�S"ML�<�#ۼ|����#��(���H�<)�MםB���5
�=bxD����G�<1�Ç�;i��aڡb`�Ց��^ܓO���u(�O�=�S¤�BHC�e �s�۟�&��)�gy"lG",*Ȼfc�7hs����)���y�Q^�H��0��#�$��y��O��z�1�
��} ���qAϬ�y(RC��U�?A���I2F��Pxb�)�Ql��\�pH�Ĩґ+��F}Ҁ�:�h��=a0�A>�R��g�*� �ȝӟp�	lX����O�N����ql �Y�b@��;D��SvA�zb2��Kߺ�
T��=D� 9`�_�#X=R�H�8����'j8D�8���_���K��X�Y�(�RT�5O�DyR�G:nJ9XC�+����W�L��~2'��O�)�Oj���>i#�\��:�b��Ǒ8���k6`�V�<�fM�iH��&k�T5P�Gi�<y��
i���uA�&/<�� �Qy�<)��8
;�9$N�Y½�eQZ�<�O�3��2&
�ڵ��QP���k���O$�9j`&15ʱp%a�m����I�h��������v�)�i	0�
�ː���3^�M��LGk+!��;m&yBQ͓�`���k��H!�d�,PD
���/�|��Aɂv%!�$
ZO�9eD�J�΍�s
B�!�$PGS.]*��;��xH�jqO��D~2o�:�?)�O	�s�  ��ڙpmr���[��R�|�����I8)a�<�7.G3@O�t[�/�Y�C�P�2��¨-��X�΅=g�B�I�x��u��
�&%^��#�
�T�vB��*H��!(9�`"E�^�hB�ɛ0��!�@��� h�BD�H2�Q�'7�-A���L"<�X�a!���C���&3���I֟P����#��� ���9�h��(�+T�B�I�-m^��qJ\�{戔s�/	�ZB�ɸT]&� �Q��\�Ї��LUXB䉌v�>���Ã6Lh8��l�p�J��D�q�'���c��ƙ��%P!�ۢ��(q�'�0�K��4�����O��[�$%h����$u��	��[�$`���&�A� � Gt�$5.]�t?F�ȓ|�@9�e�-Dy���L$A�bф�b+����`�����lr�ȓp��$0�&��i�w�>�ܴ�O� Dz��4&ɖyy�p����>'˸@
�����	��š�O��$+����m�����.��"��b�L�yRD-k:i�4O�.0E(%l��y��X���놆�
}\yQD'˒�y�g�m}�p䃏�z.*)�����y���==u��AK&q��ih GȊ��'*�#?�E����ܓ�L�hFa��]8��!�=�?AL>)�S���'(���Z#��hi,���f��MG!�	:��ѡp�Ĵ3&|���R*!�$D(7�习���@Jm:�A�Vv!�d��>�p�$ =J��9���+#�𤜠
�\+%�3y��D�G���m?\����
=��>q���^ j�`�v�Z{ج)!���?q��>� �8�G�?��L[�"�)b��""O,����s�����E�<��"O���QfFI�Ѝ��:{*�Z"O|��ä:/pCs��~����'B�<�ޯW5� S���2.�H3L�{?Q��Fe�����'N2]��`d\M�֨H�@�!qg����:D�(�GزV����j�+��E� �#D������;%���s�f�$.A�\I®!D�TK�b�+0���딡!v(I"�>D���hB��(��EƬ8�<�!u� }"�4�S��L�����J�/vJY[3D͜<�q�OiIAI�O���3������8���Y��Y� ��������y��E���[�G��jP��!Ð��y"/��x�P)X�e�H�R!�Q�yJ^��qႨ��a �1бnD,�yBeܜyd�� ��*� ��@�C��'�*#?� �Ꟑ�g�J
�pt�2��4�>l�V��?!H>��S���DX�^�XCB�Q,�$2S�]�,�!��.�B��#$Z:a�*�w���W!�d��~�U
Cd�=H��e���v�!�DM�(������E,<�Vy�Cm�F��ā+M����G^
xL"6%".��$�>����X�s�, �W�W�}��5[����?9���>I��� ��p�j�.c~��R�cGS�<��C<o�y ��w`R�+�J�<.�Qھ�Jć!�b!�*E�<�2 �gm~�`Fĝ`��;#d�\8�H����-�L�ە��> �ݡ�m�F���I����\��Y}��Y�5�آ����9��9{����yH��E(
%Q����4-�Ա��yB���J�`��)�$4RJI	����yB�[�g�X2'm&t�H8�hO;�y2�6Rzp��Ag�@بCoA:��I��HO�$�zwΚ�����$}}�=��>��֑�?y���S��q��yC��1S��Vi��C�	�N�NhT�X9T30��Q�ˣ8�bC�ɆP�ɩ�X�"`n�(�+�%tB�I���B�aҀ`
t��E�I�"B�et@�@#� ����G�U��X���<I�� cNxԙ�	J���:U�C�4���%���O>���M1��%?|8�a4�������E����s�Iy�G5�&m��[�>1�5C�D�Xu�QF�"��ȓJ8���J}R8�3D˺%����~��m�5L[�\��`6���҂�#�#<J8G���
,�(���:F�x��Rɨ�$�O0��:r=��@�շ9��Q{�M�@�!��]1 ���q�+�9`E>컕k�NK!�Ev�iP&�%Բu�a@Gb,!�_�vpi�CV=��1�i�-%��xR1� ��M�pk��<M24⃋��\�X��$�"Fx�OL��'���9L�r�&��v84��H��$�C��$q��
Ѩ�9#fԨ�j@>1C��"h��E��/לA�����%J+�B�	Lb9�ÆȀ	#8t�V"�x��C�	�q�z0�e��#�|5oZ!P��'�"=�z����2cj�Ј7�ʕ�F$�R������OH��-��	V,MQb�ɍ�3�24A��5�y��٤#�4��#w�H�jA�Ҕ�yB%A`�V%�q�Зo*���
��yb*K$���΋�R����m���yr�B���\C��#K��$C5����'�l"?�rʟ�˳��8D~�� E�MF8��O��?	K>��S��򤗗g��AB�˾`{"(��Iս3�!��  1��e@u��8���H���@"OԌ�e�^�2��KE���+����"O�Q2+_�F	f� �H�#�ܤJ�
OV�k�3+��2@@��8��e�����O��H��S+�~ ���ͼHqh��v��!+Fȵ����?	�	<t!�̇�: �A ���E�4��ȓF��dՋİt���Õ���q�����$���7(ܣ�����'�
@����+O�UQ�*�Qo���r܎- � ��I�(OD)Q�*�)>��y�5�Y>}~����O�rb�i>}�I���'\���צ�1�P��-P}R���''�e�T�;n�z��Oչcb���'c����f>w�j	����X3�1�'x�`�􇎋@.��%�8f�t	�''4� �=/z�B�.�3W�>�N�h����)&U
n(z��N<3A��IK����|�����?AL>%?��S�T��bP��N��@���?D�$�f���T�b9ص́�?U4Aa��>D�hơ��b���'#˷Q��v>D�V٘ ��) E�s���	�Z��y��Y��r㨚(g/ tȱH���'��#?�0G�ן��$DٚR+��3�Y�&��D��?�M>��S���=4.� �偙�s�0%�r�X�E�!��<A��#wA�9��h3��be!�S�c�%�%Y�v� ԩؓG-!�d.]T��4�hr�`M$���Ȼ.������-7VP�1�D�_���䑞u��>	sg-��"�u�2��!���7똰�?)����>qV��
&�(l'��#iv�r�jc�<��aA S5Z�颥�\�>��q�_�<�aP� �n@�6��$����K[�<�C�x=\H�&�P��0jN{8����dF�q��)�7G�b*����L�/����n���ϟ(�IC}-'hpZ�
(!�[*C����yBg�0�,A��R8&�H����$�y2�Еf��͛���+"P>%�!�\��y2��:�ɥ��lr�@p�ۥ�y��Y�"�����m�+Ro�� ��3��	?�HO�2��4�S:\�ҁ�&$s�4:1�>�0�ϵ�?i����S��/�ё��~\ޠp��Rw��B䉝2�8d[0΄ifzR��bM�B�	�p��a���)C�j���k�Am�C�2i��5mޡoX�Q�gŏfKdB�	4%�]H&/��IDT( !D�hJ���r���E-/��8{���#vî*T�ç!ͤj1��d>��O>�|��������pL�Vc�=�y�ȓbTȁ��N����q���T�O��#*`88soK�F-|��g�1m�,�ȓ��e.؍\�nMb!B+=L�a�rt�G���;jd�!�V��e:�=��r�D�Td�]�8<	VX+8�*\��j�/XE4���O������t}�DÐ�:z��!���M�!�$D�g�����?q�8;�-g�!�d�U��i[ �F&�ƌ"�m߬b�!��ں�Kg\;� �6Ώz��x��"ʓ{j�P�S��)��a�D�5W���E��Fx�O�B�'��Ɉ8�
B0���!�dJ��g�JC�ɪ�AH��ep���GKǋG�.C�<7<D���>�Ȱ�7!B.Y��B�	�i*���M�Rf����şz��B�	RYРs��P�P�wiɸ ���'�^#=��얶g��m9T�X�	�.��@cQ�D�7� ���O��O�OW�s$��)b�����?&��'G�P�&�"���a��,A���3��� �]ytG[�7���V��To�i�v"O4P�P!M{�h`���h_���F"O6I��*�<6���냁�E^z�`��d]�'�fX"��V���R��T�l�%���Jb�vje�'��'���Y����,J�,�@���ܖ.X����*D�� �mδ��S�Z�65�'D�@c�b�*դ�%��Mʬ*p�#D�|���A�,s�$Zu��k�֙�'�+������v���IcN:9�T��m�3XQ�$�@F0ڧH��Y�)Z�Xl���J�J���'���'�~���$j��`9�c��z�0	�'aRX��e��$��Hi��F-Y��1R�'y�Y���%}�DI U�?_h|P	�'�f�
&��F.�]9T�P�Z6�9�
�Q�Q�{��s�u���"i2re&�i�'m�Y��h���O��V\�ؐ���%R�t�>o^c4c�-~(�k��OpTR��j�g≽[т�H��F�w�� ��@��Y�v+�6.�`j�'R&�A��4�3�$�_ Y�%F8�$)Zi\�|��	y~�jҸ�?ͧ�HOL0D*�a���8bH��Ft�4"O��vH��29�g&�\2����>���i>���_}b��h`�hrV@O �zH�m^�I���
������䟀'��O�\�("mV�{�DՒ��ז2��r�N����4OP�{[��X��'�d-P��ҽWh�a��s�h��Eʟa��]��8�J$�'��	��i��?ҙz&��
L�2�m���?	��hO�c��(6�l<�|��a[9��Bi9D��4 X;��sE\���Q��`9�	��M����'k�����-`d��BW��Dӧ�V4=���'1�'��Y��!�{Q@�Y�'�<l{BJ:D�h����355�����	WB([% ,D�(B���i*lAT����iiG�/D�������L�Y��T�&3ȕ���.�� rFD=�<���`��C��1���LdQ�(��#<ڧ%�M ���]�Dmz� ���1)A�'o��'�ڕ�P�H
�x4�n�@Й
�'P���j.X�F�B
�{�@���'�b�Z�m�O��m;�I��/����'�����t���� 8�(�Ǔ_Q�D ��!\<��d�m`���Sͮ���)��|����?y�O ���h�-eڴ����L�1&"O0��Ӥ� {v�q��øq)e(�"O� �2͛1���րQ�(�4x�"O@����$GM�[��[/u�|��"Ox��e߭lh�QP.G��p("U�>QT�)�S ��M�*�h�´���=����wb/}r���z��'ɧ�'>/�J� �7=~th�O*�,��zLi��L�j�x`�u�P3�D�ȓ�0��1eӘiA���g�?�\��_��*���K�����+r>1��M�BuҦ�"R<f��clм"6܍�=���I����$�<C�!�JE}��J��"VzBL�Id�I�"|�'���vDL@�pPq���Z���K�'|X�顬�.JM�)���E�R-����'��H�B�	 P*�B�K	�BY4��	�'FŃp��3L��m�$�B�:��
�'\@@��ӻ+6�Q	A�ۡI�0�q�{�'W��9�'_�2�����7$zj�)�K>pQ ��5�'��'ߠ��2*(���lY!zc�0
�'�\k�ǖ�pL:L����wt2MB	�'R�7�Ļ5iʠ �l��}8@��'��X�_9�T�ʡ�F�!���ǓQ� ���V�����(D'�p|Ȣ�3D�����  �    �  �  *  y  �"  �(  P*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms��a?Aab��jD�O�,P���$�0y�x�����A��j�w��}�n�W�R��&R~��YBd�*���$� y�~`#_|X, ��o��L�#hZ�i$��`N:�`�O��t��XF{b� �v5��-��.s��c"ճ�~�Ƹ�R��!dH���J���7�ybf�9b��a��Ƿ��P�F&�?!D�V��|�¬�,�`sgb�i?�"�%̓@_����duP2��%�y��K%i�i�J�PLQ�ALR�>T�D��f?i�f��."�O=b@�V�DS ?G������_�h�n��0?I��Iڂ�8�L=*���ؑ�]�s�z�*5�X�L!LԢ@K��=)\9��_��0=�F�]�"�vT�YI��I!G�&\5ўԡD�U���T��*]�QHh������]�p�hQYB�G"{UlՊ7�#D��ٴ
L�K䱱"�D �2-94J�O@��@Bδ �)ۂc�T�ض�O���`ӣƠP��/0�jD��L-D�ȹĬ��s��+�G�����-��k�ڈ;��O���b�/O���'^�~(�<A'IL<{.�Y$�j��ط@Hvx��ٵD@&T�D�2��A�!,V9H��Fe�r�G���D�f��$� �`V"�q���S�˓I4�yb����l�V�Ha� �"�TA��`M���#c)��5{��!�L�����ȁ�g���ȓ�rP�5�ڛEC��!dO�	&���	%}(�X6 @b��a��Y�;���)��40V�e
�Rw|��&�C������4�|���62�V�h�����8@q�'`���I.�5��é|�D�ۺ��'�J�(���j���ɕ	��s:}@�S^�}Aw�ܟ2ܠ���� 9�
7n4N?���		P�8	����P�v@��l��VCY�-��Q��[n E{ @@6�QTbóX�4� �Ɇ�~2�J,")��"@a�"� IZ!L�-�y�	]5'�ҝ@��(�Ҽ��"���?q�(�$^����*Ż(l(��Ue?�r�K�}`k1��Pd(��f#��y��{�ir4�
hjR\���=���5
�v?Q���f��O��@Q�$��@��r&�d�f�#���1�}"���$q�Ț� �����G)~��%*������H�_HΌq���(z�bi�C�'��4" ��k��)�(����EI��$��͈Ȳ�Œ8'%
%K2#4U���0k2�� ���������O�]f!� �a|���W�;M،i[��IW�#�^% �҆ɐ��J��v���~���IXFr�8�Q�)?
@��l�E\!�dٛ'i�*�KCRi:���ͶZa�x��S��~��f(6�)��ii@.%�I�{8�ԏL�$�����2)B��"!i�d�����Ed��°��Y��1�0�+T
�YFB�=,�~����)�n����3�Б���I3j��rd�6ў,��*T$n�hЈ�!]� �6����ȓ$�Z��� bBE�&��d���$D��7=:N�X��M3��J�i�	��̞^4�2P��6�´���S�'QƀRp��;R���P'F)H�.!��'��4���R01�g� xt|�8�*G��x�#����o�Y��gQ1O�٪D��:R\��f�/V��4�""O�b�@�TY6�G/\�]� ��"O:P��F��'j1���20���"OR��!�CY:��-ƆO}�<`V"O�����+]�Yr�͝�]�5;`"O��C��,���R!�*v4�@"O���e����4���|V�\ۤ"O�P�#/I.��zU�y@�M�G"O��iҎef`�b��z�41ia"OL�P��
eڰ�B��>h�Hȡ"O<����&�&,�Co��`�����"O�aQ�ٮAf���ݞA�a��"Opy����L#��1BM�4%�U#"O�,�l�>p���$/^IwbA�c"O��؅��&Q�H�aM�>?�dr"O,aYgi'A-��BR�:=���Qg"O�����gH���S"ۼ#�H�5"O��@�#S��I�D�23��_�<�MG�:�m ��/x`�hq��W�<��hڜ&�|�3����"@p�"V�<!�o�?l��aV`��a�j�ծ�Q�<�uG�\W ��𩛔mY�iNTQ�<��l k�8u���֐<��%y�e�c�<A��DIU���'�s
ԡ#$JX�<���<�
�H�I�X��a��o�<��\�-7�!���>Uɀy��C�<�ŊҞ10h��> ��Z�j]�<'�H��z}�Ì%�� t�M�<Qe�9��@`r��5<xt؆"CH�<�QW9<ī�-�n)�Īs��\�<)r�Q��,K�� +���
3E�V�<1s�=f\�zu�7�Ig��m�<�uF/��|�4k�+22n�t�b�<�pbV�D���I�Dg��|;A�a�<�W��3��s�	�t��}ZG��h�<q��ƌ65.x���k��5r��K�<)s�
	�j���zP`C�<��h !�4Kfj,i5��ˡ�@_�<��;yFy�dϩ�l����S�<YÈPV%Y�@ͼg~9��OS�<�5BZ/Bf��{��Գq#�!���CQ�<I�i��9�X= �)B�z@0��Y�<p/D�'"ȍ'�%��cU�<�4��#m8d���K�jn:<{�I�<ɧ�
T	|}Х(īL��0�A�D�<Y�j9�p��q!��ܹ8R��h�<�q�W
��:��$^�ʙ�EF�a�<��e�,gV�l�����\XȔ��B�<1��ڦ"�䛱�ײ��=�Z��ȓ<��(�Ǧ��*<��.)a��E�ȓ-
�CF ѳ5a�c�Ο?q�����S�? ��@BC��B�a��c��h�"X�"O�a����4�@K�B���}��"O8�ā^!Of>p�3�C t 9Hp"O��G*B�zD�4!��$BY��"Op��A #+:�� ���$._�D�"O�9����8�Q�M�DE��j�'��*H�9�4�fEE�_�6P��'U��8D!WQ�\HQ�^nU+�'���1`��	h,㰭�Y��Ls	�'����͂�mϲd@@$C�V��r�'8��ʃ�ޒ;e���$�EO�>��'Q�H&d��b{�0�T�p˄�	�'s�PC�-!Nv�h���}�Y	�'��};'�@؅ic慭t�� ��'���s#�G���k�c,i��0��'�Nx�" O69J|��iׯn�^�K�'�l�z4�R�2L��` BH�pN0�'!:̩s ߷r
��3@�"|ծ|p�'Gmh��6�^�B#�x*�x�'�+o�61h (%�.!�U�V�/D�` f��L��0��8T�Y  N:D���� ԛH9��{� ݔ�����&D���M�mJP8�癢k���R��%D�t�%!Y�,@�i�v�X�9ž�Zc#D��V��Q0����o��P2�<k�d D�� S�@G�����Ֆ.^yȆM.D��A+�9Æ8��F$�>��`�&D���5̏�u[̑�Fj&2[4A$D�D'���+J��p��#g�2�1!-8D��+A�יఽ�T��_�m`�1D�|�t�;;8.<KAM��ۅ1D��p�B��JΊ���",)�<�e4D�|�*V�Ghn	�R� V�t|��(D�h�T�\��8R$����K�f5D�x*HѰp�u�@�b���W` D�j#���>p�C�D�|8���"D��� �I�q�M��Gn"<q��!D�4b�)ރ�f!���P2���j@m/D�4�P�Y�Q"P�2�O�!?,,��7D�t�J�!>T^+V��5T`�i�6D�<É�/�nhhuD�#B"��F�2D���I>���S3IC�	��4J��5D�<+��1i&�ɡ&l �L���E3D�tᦨ	{�``2
ϯ`?|�!"�1D��xR�^�����O���"s�?D���!!��m$�I�ɉn��B6�!D�`('�M�N��p#d����M�W�,T�pr�*�@����2hֺuؕ"OVaʰ��t�`��p
��=`"O(��LP$aVV�q��<]��"O�aJU�[�?�=��L֋xYv�bR"O����*,�,@��V�
_J��"O�x��k�X���"�l�n�Hq"O����+��"��vȶ�Pq"O���O�%��ՑD74�|9�"O0���x/)��O�2���J"O��c�m�ϢAc �H7'�2� "Or�y�̘�{NѨe&םUBB�k�"O|�
��%0�2� %	&@ȑ�"O���𩇡 G.<�&���t�"Oq@�I�l�\ �B��r���#"O�<�7�ɞm/ؘ�oƱP�%x"OH)H���@�Ne9.��sz����"OĔ� �ק�r�{�NS�Fx��&"O� �X��N�C�j��5��vq>��P"O��a]�- ��kN
*prmi5"O��f�/�X�	���2F�u:�"O�Ih��B<&�
��6`<ƒ�k�"O �r�Ā(�5��-T�G&��W"Oz0���ә/"l�L 3�Ģ"O�8v�s�NԺ��:����"O�A�&^�81h��t�ڏ��$�A"O�A��dY������GͰTy.�֎{���/B_X��J��!h�؀i�̋ ;���@�=D���I��xz$��:p����<D�HL��X����ؘ��=D�4�hC/VD�(��׾�\����1D���c�*����
	�N�[�,1D�p�T�N���l�e���Z�,,�e`2D��@�J�q��(`!+�z�<�&�1D��P��w��XD�.��0��*D�H�
��q -H%��I��;��)D���g� �?ab�i@E�S��}I�,(D�L��	�_��9�6#
��:D��)��˱H�Hd���D�RJ�S�'7D�S��=6Y���E>aT��'F!D�x"��ѐ�j�zjN�M�X��� D�3��A�z�$��%@�8���+0�1D����ջ:ڢ�B��wv�]�� 2D���	g	Ƒ�wj�1�#%%D���b`F�gyn$�fǋ�q�~	��I8D���T?���4(=�����8D�1�%U�{o���*�C�f�X"D�<�%2BW��"M ���K"D���eN�']*mBC�ðSx&��!�"D�<��X=Lu�d�򩀼-�"x �@!D�T��Hߺ�HT蜔W{4dB3+$D�����={�Y�"�P����!D� �r�¤��K&g�q4�a;SO#D�0�2�^����ĭX����ej%D�t�c�F�<*4�&�@��׉!�$��(>l�2�T�<[bI�.�!�ć(hЄj�-�t �S�!���[��y U���`��M�@!!��!#Lv�P�ǒ���D�c!�Č�J|8��_7����:{�!�䈸�h��򎊴 ?8\�[>�!�]+�:1"Q�I|%��*�+\1!��M�U��JE}	h;Eܭn!�Đ��x���~�B��E�Q!�$�_u>9��A'�H �&��!�DL�,Hi��f
�~ɨ��U��!�d]�����N	~ D ��%v!���������3^�L�Bp�	d!��-�}�ģƪR	��Y�J*D!��ҺsY�H:�'�
S�@��e�,V�!򤎿b��� B)C-�QY�D^%N�!�d��GG�p6�ͷ>�!�5^6wy!�M�-P�G�0k���4D�c!�D:/t�Ȱ�)�]�@U�c��S�!�	'�T���Ȱf��DI����#�!���}�$�2�"�t�`̹��1	l!�Ǜ.������ծC*�j$�\j!�#�$���n�q�*�qFe!�!�ēq�"���'��v�L,_�!�ǣy�$A��DK�X���fd�6�!�D��5h�q9�LY9i�m���Z�mN!򤐖q(�����c��	
"S2!�� ��YC%N�o�Ha$�_��-Z�"O
m�ǩr����cA,lF$�V"Ou� ��T�
��ͼB+�Q��"O8S�a�HoFMA'FF�$�<��"Ol<!��[4H� �g�'|g�|�G"O��qA�hS8g r@E��"O�`��F`��81����:;�M�e"O�y2kӜ%y�,�����u�S�y�L��0!v��-�,�xt�K(�y2�F$E��qeO%#�m��,S�yr'�)dH1���I�$�h�� �y�ĝ�*9�y���mn�Kw�Z �y�n�
s~Cbd�"j|X:N��y~"����
^t�=j���"�y�"\�������[�h��˻�yb�L�k<ܤ)��N!U�H�f��0�y"DՍ>�D���Z�i��4��N��y��*ֲ�r�j�b���� ���yR��0�p���m\7G�t��)	��y����44����ד��X��mP5�y"�R�
�ڡhӄ	z�24s���y�oY8NJ�aǠQ�_N��j�7�yB�˭7~)�Ώ
w(�����y�K�ml�@��L�Jxu���y2DT�%v�!����i+.�y2��>��Â��z�����H��ye	/l�t�D(F%$)��ē��y�,�aH5(4eJ"xp!Cgπ/�y�)�Vvx�n���8�q�[e�<YaD]!5�СG��eQ[��z�<)ƍ_$1x�]%�PL����Hs�<��`�*��Bg@?Y�S��g�<A���cĸa���)z�J�de�<Y�*��26D��N-5�P1F�Yf�<I����Vd�Q,C7����&l�<��͊X�@�q�P�;�,sÉFk�<����C�t�2䞅~�)K⢛�<��/@�R��|����LdB�*�*�f�<�!嗍i�L�Q����Y Ѣ�dZz�<Iqi%v�*T �K�8�r��Nt�<�s�QY�����/"2Mra��w�<��%�0S4�jf�0Ht�Bc��]�<�TŃ�[;TTA�Z�7_�i��i�r�<AB��5q��i��g\-K.n ���j�<�U����y���ڏ\��2#�M�<� m4���cM�Y/TAb��J�<)���/	z���F�'t�>����G�<9$�Ƃ�ph�#Q=��Έh�<oR�}1��镎�D/�I�Bmo�<���b�b�B[ .t샧f�k�<�&Nƴh`���"p�$��m�N�<A$�	�:��R�	C�]��� ��S�<9���2&ּ��k�>f ����a�t�<�@JVj-���!��j��(�U,LU�<���?���!�Ο3u ��w�CQ�<QF�Y0��`�O�tl�"��M�<����?Ճ��N���s���J�<�c��$�j�Y��;)�� 3�@�<B���q�y�VMA�6���"W�x�<��ME�'�j�뀮�0h.Hԛ��v�<Yr��r�D!�#�,J����g�<Q���)��4��l��Q��{���w�<u4
��ib�ʇ�72Z Qb��r�<Q�'P Y~`�&H>'r ���,v�<� 
(	�GɈe����M/T�ӥ"O<���CF7,��
�6\��A�"O��a�NS8V�j�s�H��/� �"O|j��"�%�?D'x�yc�A��y"m�L�X��4Rv2�dY5�y����� �`�)Lš�-��y�䍘��艕E��Q�tY$+��y��է=זѲR�L8:�p`�ā��y"'�.)&����9�`A��`X��yr	�<0�J�QC74�Hg���yb��ZLɸ�8)j�#�M��yr��C�8��c����9&#�$�y�@� ���m&�6��I]&�y�B
CE�I���M����k��ɟ�yr�X��	��*P���V��yB�I<B#�)��D�>U�n8V� ��yJ0� �86&ݶ~1��h����y���=äI(���oJą!Վ���y�#N�#��/Ċ`:���f@
�y�)�9U9�s�T�QHErD��y�o�>�4Ht����P��D�y���8M�5cnB et �H��y����
x(cAK����F��<�y�JK�,�B�˵�+���S+�y�IC�:m�[��ҫ �j�9�,� �y�D f�%�C��x��$�3(�
�yR+��	�	���O�h1�廇�T�y2B�T�\-��	ozT1�J�9�yB���Sj҄
eH�{�l=������y���5y.�A�u�΅c��%X���y���"
���1��Tm�FEc�$�'�y�	�>�x(P�OY�c�f��@"���y�߶[plْ� ��u9����yR)&?8�䙑��X��1�r ��y ��`��iK��M���1	��yb?�P�8p@�v6 	��)���y�`C$P�)Т/4�ZH���y"���'�<�襎Pc������y�ݙ��Q,U��A�#���\��F>l�Q�]�o�� �n׻�FĆ�#ڞ�˴%�Uk*�k��l�(��R�=���׆>p����H�%���ȓ$���+7�}�A+p ɐ�����%���>k�T(���^.�*q���jM	��ٚ 5��A�+-{����+����@�fYD��	�%'n渆ȓ1��ņ�(��h�I������)z����P@�#fD�<���ȓ7$���>z���0�Ɲ A� �ȓN@����M�'�6�C����$�te�ȓ�D+�L˓��\�D�V�4��ȓ0�hx#0��,QN\�'J��&�N���ҺRF�
^F��9mH<��5�H=(qcA�,���&Y��l��|����#�W��т��O/U��ل�E*Չ��N "��XB��èC@ P��o�6�aP肍Z���1�	I" ��-��}`���QiA�d^R ����t��i=0�
GaI>yLl��E�ʘ	(d��R�Iۧ#�.�U������ȓ�~�۷�^0z�m�Q�F±�ȓ^z���"I�q���c0d��Y��ȓ��@A��Ch;aJ�5�؇�l�|�@�(���W�G���m��S�? �T�W�G�2m�p�K\�vp�R"O��Ô��*?4�<r%��
�x8�"O��SRk��
.A�Af
�M��i"O�,��_M�vL[d�M�PQZX[#"O~�򢏂	X�(8��ċ=o4Yj�"O��P����B����3Ȍh�"O�<�Ǥ�	�F �գ=�N��"OTM�ğ�>\�1y��Z	�,�"Ob,�ҁKZd� ��@�2>}h ��"O���f���<��
۝OxUp�"OD�fm�v�F�����e�� �"O�}� %�6,a��3[RV-9e"O�(�F���{��(� �J�ɲ�"O ��`�  ��   �	  �  �  �  B&  /  �9  �D  �O  |Z  de  \p  /|  Ƈ  ܒ  ��  ��  M�  ֲ  ��  1�  ��  +�  n�  ��  ��  ?�  ��  ��  �  ]  �  � � i   ' �- �3 : T@ �F �L "S �Y �` �f Jp �x # g� � �� � 5� L� �  x�y�C˸��%�RO5d��pJ�'l��I�By��@0�'�F��A��|�^{���OM4ؐ�Їv�lh��Y�&7�C1Jɜ��AP�Hj�%+5#]/AT֝�ҍ�"�x�S(#�t�	0�� �Pp�h�� ���rI�	cUhm���>>O�|�6k�p��`Xw��dU�O������q �P4b�d��A��$lkL`����t
��Ia���9A)�9��=n�<;� �I۟P�I���ɘ(ɼ4��M7P(� �c<w���	���I�x�'���t��ϟ$�`J�4j� ���~���eFşx�	J��ß�ɵO2�y" �l/>�(fLѓXi�q�Wf��y��+N0�*�XҮ t���?I�[�qV��q�՟>0�����uH5�Q�]:ʙ�襟8�@dܚ#�()`�ҵ�,�B��O��D�O<���O����O���1�S!O2�A��>b��'h�/6������������'E6�@ڦ�޴!��	�1�Q�V��9q��w���b�ԭE{��O��=ke'ԥbhE��P�o9Aϓ�OT����f�9���������G�'wў"~z#m(@d9+�nQ��"��u�è��-�O`@����]w��"6c��M����[y��p�Ҽ1����2��W��8c���)�n���3	���B`�I�OѴ�����:�	�>���@�QS�.+g��Rte�'Jt��9�D�Ob�?�'+zI�7��4���:A�Kx��!�'�By�ЭB�XE��,��u��+�',��k��0��I�m1ܩ��'rʔ��b1{W�^������B4]<�}ȳ�Q�l���7����hO�U{���.;�  X��"
��	�$A���m�	؟`���)�y���PtFi�/�1*">C��g*@�I���}Uȡ:��I0	�(C�I�d� �*��Y� ��M�r�ȭ�JB�Ir>��!w�Կ:0@����J�V�?)1�S�c��jshޘuZ<L�S�Z���Ix������	c~��{�r=��eY�� �$��y��˅"ب-�`y2�,��mI��yB�:_���kR/I�n$(�r�GG��yb V�"C<$R��G��h���y��E�=�hY��
�����d+��
P��(���1��3B���1vz$��S�lp��ǟX��K�)��60��қXQfY[c�˳+�VB�=`߼ �%�S�>�M
�q��B�	�?��[E#��'z�p�u�ɿ{�C�	qR*��4l
b�`H2È�@�rC�'7���(5 ҙ?~���DҠQD�O^H�>Q��U�<��O��9E�9KQ����/�.C邕���'��'��6��1�7��� O���T-T7*V"��Qi<J㚝��A*O��1�cd>�;L�,X�@#od�5�rLߔE����*O}#��'�r�'W`��D{ȸ�V(N<;$
4?�I�X�?E�4A@�O�pE0��/ ��XB� W���?A��'�6 �� }���M�,/�Mj����d�;:���$)�s�0�'@�P2��R�vk�!�����=��!�	��t{��/�|�"|2qI�#>�f��h϶US��Ӗm�D~"cX�l��=E��E[
�`��	A�[��8��Z������@���'��O�1��Q�E��1/R$%��
�' h0��|��'0az,�V/�A�t	�*{�dyr��O�@G��h �*w���&'J�p�H��?Y�(�3��'T�4�'.╟�"A��f�(��2d���҈cM9D�dcu�P��x34��2�X���$D�LS@��M�^�:ԫ0�h��=D�p�Ňhܘ���T-z�|X��'D�� bl���֡T�
�`Dꗈ�<�1�)�'r^���J�-�$�.�%��0��j�<����?����S��ݡ�<C��1G8@&|�.)i7O���`�׊R00��IW�ܸq	͊J|!�䗊4؄���F��MR�c�6��P���'l�'=BX��g�62Й�C�\� w���q��K��
�'+��˕��!��;a�I�G�VM�I>���i��S�\��O�j�Xa�+3����DV"o���	H�	��'6�!Gx
� N��o�!5��4S��
�V�����'��Џ��	�X�䅐�I�k�&�S��Ǎ4paxR���?��y���	���5���ʬ�����y��g*. r�I��",2&a����?A��'�D���6Pir�H@�8^i\�*��d��nA���(W���Ǫ�5�< �*ӥ$���Iɟ��ɽU�t R"�"��gk�r��B�qT��5�W 8B�}����/��B��9%�s�ݠ2S�ѻ��T�K��C�I�wĵ�%BB�B)di�@� V\ޣ?� 퓍h�)�� ع�b��!+ߖ3X��NS����D�Iz~򏒟,e��'�L���������y����5�T�B�v,�"�y���R>��A�!RZ�!�f��;�y��Tkj�!��<�8؅�=�y�,�-_��S1C�42�%��P���s��(�7��i��p($(�-Z��(PZ��h4N�����Im�)�S��.M�G����".Si�kI3D��Q�F�P$�a��њe`x��F4D���%#Ю��И��.
�~q���0D�� ��
�1l�thwb�=@Ht��F�.D��� ��w�@�x@Oį d�Q�L.��P�'MU��'
�A���w�C��]�������?ɍ�L��JfQ�)��x��bV0p�`�*��!D�8:#i�!j��)0��Ӻq �a%D��b��-.�b�卆z 5 &.D���)M�j�Rq0��.������-�O$��Ig7��+�7��s��_PƢ=��)r�OT�X�F��B�t�� �O޺��'4B�'�F���(\�R��š�a�z�'�y��U),*p�KSq����'Q�P%coz���銫DNr)��'��|!f�R�i�L�S-��-��
��dGb�O�j,�p��:tDɁ����P{�u���Ex�Ot�'��-"d���%��R�6L�%D�B䉔�+*׆L0������!8v���'y荺a�c��y�e� ��u�'�T�r�`�Sd��u,�u�Y �'�x�)�N�W�δrga�p�$+O�0Dz��T&,IL����� }�F����5"c�99�
��I��%��>u�â��X8�{sk�X{��3b�*D�li�I��Ut�����3*Ȅ�h)D�,S��/qÄ	���[9����<D���'�$��r�O�}���&D��T�;���S�KH����&>���r�'�:���' �@A�צ���:���&'{jqb���䓧?a��L�\3�ޮd�z���ET�=�d�{q0D������0^�'��Br���/D���	�Q�`)�QcLr�4��,D�PqAψ!8�I���8���P�e(�Ox��I�ls$%�R)��N������0q<��=���c�O���c'��=H�Z�bK�|T^-���'b��'�jx+��C4\��[����
�	�'QP�;�A�5��x�%*�
�b�	�'�$��E��t�t`fC� N�N0��'
�A���r�@y�֡-M.����d�~�Oo08FC\�0��Q�v��"K�����:(Fx�O`B�'����C��	;��v)n��e�!_�C�	�P<�R�X�DǤ���*�;,rC��&��0g�ˁ}j�s% ={nC�	�t��X#E�#M�9���$:��B�I�h`���ľW�TYG�Z�mG�ʓl���|�Q�f"�<yN�#a�DP;�LUyʇ6�B�'Dɧ�OK4��G��`ʨd٢­d�40��� @��D%S6%9�)RE�2S �P�"O|E�3��&��`�����C��	"On�V�I�/Y��ң��b�|z�"O�� q|�92�kN#K��`࠙|�1��΍�W�E����e%`mx�K��~Q�I`�	�����ON�R l/��i$�^1v� ��V"O��nV�H	�r�ۃ�$��"O����� `6�iӳGU!xᆌ"5"OL�30ʑ>��|qQ��&b��,ٶ�'Բ��Γ&C�Q1��c�DxR��&�ўLIK6�'!�ݨr�ؖN���Da�5^q$	C���?i�j�lx1����V ���a/׭%�D��1����ͩ�jȃ7&�'m�m���0Eq(�V	�Tc�fR� l:�ȓb�d9�'O�/$zx+���j:�D� ڧ�$Icf�6n�0�+G��,�F}��-K��"<�'�?����D�"*&<�7� ���!�ƞ7!��J2b��w����Nh0�G�I!�>0Ȉ�҇� eR�,b�`B�u*!�dH*�"��Iţa���DJ�6�!�d3`�$ٓ��t��ъb��{�剽�HOQ>�'�<!�X��dg�C��U�BA�<��M"�?����Sܧ9|Ѡ�\�0��M0�eƪP���ȓTp����r|�X�2�C>U��X��@�n1Au&V9���J�9��t�ȓH�p]��G��j��� �L	5P��$���.aY��lV��
����$�D0��$�71<�$G"~P���F�k�^���H�.�|��'N��Oծ1��5V�,�F')
I�ȓ+;�4�*���r؁�l������).>��G��@�f�:��(���XL�G	De�8�P-�;<=�Q��Ɋ�?iƉ��kX.��Vhڔy���a�Xt�'.d�َ��N2��!�uJ)ق𰫉�-/����O��d�/7b2��%g�]&�0���<c!�䇗=Cd�:D� %�`Q��u\!�d�!���
�&
B����0@L6hR!�˹;��ŀ��Ph�,T��?">џ������2G>ܨk���,�����<< ,R�O���O���-?�A���=-)���0P�b�D_�<Y��s�`��%�[g��!E�Z�<9�I=�tX�G�k գV��W�<c$S5�
�� E��eF���Y�RB䉪(�nE�󣊺�PX�#� �U���|��LZ�A,������ ��K�Sy�c	��'^ɧ�OY�Pk��!x~����ʗW��-�	�'~��ir�Ӭ�\E)`�PDd�b�'p�X)1�֠�ݣBO|N̽�'>zUC���cY��1�Z�%�b���'�H�cE쒛U5�m�6%V�2�܁�M>����">��t0<q�EK�zĀD����45���1���OB�?�''�����j��j��H�C�(K	�'s�	�S[�,;F�V&@1l ��'��8�sf�8
~$��iG�A�4�	�'����A�"Ore�׀c�6��� Y�U�fPc*X�CdU`��E2�hO����Ӫ<زS �hvD*'��'vcxD��韐���6�䲗G�5A��I�#Z+vB�	>�=���2i�t��냜n�B�ɶ`W�`	A�H*z�ah��*2.B�I�Z����I���@�b�
!ܢ?A�5m`��$��'UV͊s/��Y����"2���S��,�Ib~B��N��k��]�\�R͠DCִ�yB+�6%�dy�&	
�,���+X2�y
� ��	�.΀y��o�Ը�xf"O8T�Ц�1g�*�x�0]T�
@"Ot	�n\�ȉ��)dZ>���Q�����哮\�%��<Pe�g�]#}�0ʓd��R��?AH>�}*�I��*9�0�n�b�����
�]�<�5C�v.�j`�ę%��mc���X�<���(z�=ku�?8��m�%M�U�<�L�bP�\���6+)�؋%M^M�<��
;F�E��
�W3 �h���d��1��O�� ��OȌ�G�G����)�������'�'���>��GO
e�������t�4�RWkKQ�<�!C<`����%�ȑ5�۱�V�<ё��j%z9�6��X8��U�<�%"E�'�%I�)� �~���C�Q���R�b�ȼI�/��1"�&�D���D{l�͈�܄bFоhϸѡ���t��1se�O���9�O�I+�F���@׮D��"O\x�rF���0%�sgM�H<p�"OH\ȰA��p!���s䌲y'�yc�"O��ٔ�� iiT$ #�.�<(�g��%�h�|�	1�Z�3�<�8�Ʃk�x�$�'�Rh���4�H��O@�)�Ո�B9$l���?�~\�ȓ4�z���V��B�[e�Q_����kP�}����$LAJ�;�aJ��d��o>��p���K������Zذ��G��5�Gn�*�<٪w��|Ӵa�'T�#=E�Tb͍_��Y@���i���J������ƈ���$�OƒOq�<��sƁJ"�� �O%{�<b�"O�U����J��AK�,�t�p"Od 1����L�2��c�Ɲ'�>�*�"O�X@ƛg=
���n�(���"ORs�ٵY����Eڿ$tX�(�|��%�ES�i�9�4��'�!*4;!g�W��(��e�П���O$hp2� �7�<��+�;V9B�"O$!�E�ՁZ���S�TIX�Ӱ"O����bO%���1j��:ij �"OԸ�G٥JaHвh�F^�M�f�'y*�$n�ܰEί5��@3�$Dvў$r�O$�Z$^�	4�ʀ/ƐZ�"Mm������?y
�M�$�M	u�dP��T�[�&Ԇ�9~B�B7��_��Q2�ȇy�Ȇ�I��AQ �37��L�w��Vt��ȓ1Ŋ����Ak/��p�O�-��HF2�-�'![l	Cw��g ��T;����I�H�"<ͧ�?�����AM Dz�&�#[�����m��X!�d�3p.~Ic��_?C�̭��k�`�!�$K*I
P��$×6¸���a�,�!�d�	�Z�@�B�+,�*ڒ��9%�!�� s�Ԙ��+ �X�����<�創�HOQ>%���S:K��s7�/M=H��<��#��?!����S�'z�ހ���)\I!mͺNu�]��Eb����h�G��P��&_�^�͆�DD�)�b�ԉi�Fe
L��[3vy�ȓ=���H��ڃe�0b�D̙��d�<�!'R��t���B�:�d��g�g�:��O�#D�O�$B䉥���2m�"�&���'Q�'���>Q�
ӹa��S�0Z��-�`�i�<��L�>=�p`���R�B���e�<���=gj�1��M$n�D!K�B�^�<!��1�~� �G�t�D3KR�����f������ (�nzBȒ#~�E{�kF�҈�Rqq��Y�b/x�H��IH�y���OX��5�O��b@�͘�3�ڗ
5�h��"OFD��ɓ	"<�A[ �`�)�"O� @�8fIP��h�rr�H�0EY�"O���p��m��H���`����	��h��B�M�n�c�ʚ�6����' &IJ��4���$�O��3�V`�nLq�&2���f��=�ȓ��1£Q2M}8Tae��*(��ȓ=�L	��iÚN.�$�Q���Ԇ�0���E_�pIH�
��V5���uz �2L�f�K7O-�$�'5�"=E�Th�M��lX�iB�l���Zb
����v��d�Of�Oq���S�A�Ct��	��O�o<N	s�"O�q��@�(�Jj�4�J�"O�p�"ءiu���ɘ.V8Ȉ�"O�2k�2Y�� +،~�HXf"Ot�SF��	�f!2c��N�
ĩF�|�,*������M�c�;�f�鰅U�T�L��@�	�����O<x#��&aY�ɢ�E	�)r�8��"O�p�%N�w�2�TNNcS�a)&"O*�Av���E���c�Y�O7�h1`"O��#��0G
2qp'I�C?���c�'Yh��Յ-tbhҵ��(c��	
 ��(�ўЉ��4�:8����X�Xk��W�t�����?�t`�X�ă?"�ڭC��]+YB�ȓA����MR�~�
<�'j�*g��؇ȓ_�8�S��ݫ�r9�'�	�{WJчȓƖ]׌��"�,Dσ�
dr�E��#�'c�60�H�0����@�S�°���q�#<ͧ�?9�����^<U��TBSj��T���� lN�u�!�� 	���vmD�g_ؠ��+�22�!���Uo�P�ǫ�U.P "� ��a�!���2*�`��ǌ1���`gI�!W�!��͌]BxӇ@
4�VX!���剠�HO>}�WՑx�� ���)r��]��nY֟�O��'{� I�O��'���RU��&h�^�@Fꖫw%�����|R�'E��4o\fу',	@��	3���O�!1ub���KWx@=S&�z8��Hg���(a�C�Q#��Ozt pB�d��š@�Ȧ����� ��'&1�R��uK�H�4�j��[�U���pR�����=+�ӆd�:6��ab!&��	�(���OLyr��	M.�b��T&n�hUr3#����D�7Z����O��?�	���� �/����2c�"���Aޟ0
O�Hp��,��Ku�X��S�O)�HeG�, �5�&#􌩜'&*Ѩc�l�Z@�"Ă�}N�?-���׷p�Lia�	"W#\�(6�s�`S '�O���#?%?��'p�hI�*ʿ��a��[�4J�@	�'Hz��$�*6�\�y��ܸ���1��$�m�O���R$LK+jr�(�f�!��V.D�:��O4�i�O��/�Dۍ2�bL*��[	ˈ�y�IO��B�(vb^БF��	?�f];�
��ܜB��*S`<h���2Z�8��wE��]_�B���đ���N1���T�&=~B��&[��C�M�>�y`��T�G����B�����H�`��62�؅O�d]F-�U��O,���O�d6��ӹUWh��"I��K���YR;Y�~B�	�`��Li⌙�9�`� *��.h^B��	-�H�	j4=��X�2B�I�
�����* )]$)B�ɫ,^�B�	>��c���\Z��G%/;˓`ӑ��BC�6}�@�;/K��p�f�9pX�g#�'�䓓?��0<i`ߍe��� �q���A���S�<i��	Ǫ�6�f�hDO�<	C�BAQ&$+�O >aЍZ�-b�<�,�U� a���`��|
0d
ax���/O@�X��F�IT(pmާ!�f�8 ���o��������n٫,:�����u���������� �f�("CL�L��!CG�}:0,�ȓtҸE��� 	�8D�UX�l�,4��S�? �eHchwѼM�dbS<_r�U"O�Iٓ�CJ�Z�i�&^�C���蟆,�J1�t\���.e{l����=�O��)�O
�$ �56ȑ�sg��x�V�X�A��6�zB�	*\�]z�BAg��(5���TB��
�^���d����Т ��qm,B�I��\�!!UQɞ!���%v\C䉥B��Y2�!�J��	y���vj��dCZ�������oT,�^�*�B�1i�cA�O��:���O���,��5LL:�r��}���F �sLvB�I�"���RBM��#��NDC�Ɂ4Vm��5��ج?~:���o��|{����R�ƥ���<W�t��ȓN��T��C�0[+@y��%�5
`���'<�"?	Ӧ�g���,�������H�b$��ꓧg>�'���'.axB�T`zl�����^��pӲ��4�y����0ǎ��KƳWD�"�ۍ�yR �����P�KN|����n��y�j<Rf�a���K����E���$ry���i��1�G��J��3�@W����O&��<���kz��3����l����)V����O��xKB��>�©S����;8�@q�!�����&�d����|B�NЗz,!�4�W�4��ɠ�~��W;���|�t�l��R+ �(h�E"P90�0��󢝣���DD�d��KR�F�O��$2�n.��I3	ˍ8�`Q����]��RB?ٌ�9OR5�5�6n2X{�їg7b��e2[��-��"�PD�O���On�I$�Q�^Δ�j�.�a;��F��O4,�v�S"u�>=�]���"p �V��8�	�:�.�'��'xHآO����4J��� �Nז�
�KN�];�a�'6,]�I�x
���٨^ �aRG�2U�V����W�3��5��,̔U�O�s�X:�+>?	@��p�N�t��>��ٻ��AV�/O�HW���3�ӲB`�E�%&�?
'���ܘMP"�Dۇ�~RF�(���?�	:6����2���zD��+��@h"����'lba��	h�����*��=<)2#�1_��B�Ɏc���ᢍL���}Ba+
?@�B�$^Eڍ���Z�"��%�2/�r��B�	�s�`���ՅT��Y2D,%fB�I�~;����i����27eBB�	C���̝�yN�;Ӥ �cB䉸qU����N*@v(k i_	PC��,A�R-:d���J��ɖb9�C�I��й�MZ;.B����nC��L��(�� �v�>�P�$ԥp-C�I�e�
@+f+\/�t�тc�[��B��?'��]�LΖoJ�M��ĲR7�B�I�O&��+5&�% �9��8lX�B䉍��lJ�)]/W^� Â���!��#?����?���?!�[p e�� �c���<W��)�i�b�'Z��'>�')r�'f��'�0��֣&���aƥO(jغ��e���d�O����Od���Oh���O,���O����̟|�6��3!&m��X���¦���ǟ8�I۟X�	ܟ��ğ�������#��l0n�AS�
>�d�K��ז�M����?y���?��?���?!���?	��ZI�X���ϦJO8���0����'�"�'��'�r�'���'~2��8���ps�^8(~�	3PB��G��6-�OD�$�O@���O����O��d�O��dY�B����ʲf~i��_"9!BAn���H�	�����Iӟ�������	�0���ٱO�#Ӿ�H�	��?�~|��4�?1��?Y��?i���?y��?	�E;��nbԍ��K{N���ÿi��'v2�'lr�'���'���'��ഩ�B�zL�Db�	Jzp�
u�j� ���OF���O8���O���O��$�OT�Aw'ٴy�<�Ec�_C@��`l����	˟��I͟|��ڟ������	�i@fH�B��4�Jb#հ;xt��ٴ�?���?1���?!���?����?��qZ��t��]xμ�����3��i\�I��'?Ib�̘�CA����P�f��D�6
o}�T�\��D�'�?�'LZ���e],M�J`,A����s+R֟h���<��O2��L�8#�'���ÝA���K$�w���-�28O�e��.X�ў���<lǿs���I�������'e�'��c?��	|�? ��UjФ)� �r8/�L��"��<)���?�'$�.>0dQ�B�N�U29:�ڹu!(ʓ�?�e	�h��1���ҟ�cR1O�l*�n���V�B�
5c�Q0Q���'b"��:&�  ��d�g�:K���c��O���'��I�p�?�'ڸ��v�^�����2�D���?i���?���_5�M��Ov�Ӆ��^w(�\0���0"�TJL�"�A�����ON���O����,oe�5`�m>�0R�<�rY�x�'���	��6^͊D+]�dp�A���Q�.��ʓ�?����yB��h����i��8�<x��E�"a�oܠn����?�p�O8�I>�(OD�[v��3�V1��ҕM�l�4|O���'���y��ʒ����=G�"�'��Oʓ�?A��y��{c*���S�����%�:�)��4��$��i�֘S��O�"�����ݙ.�ּE��=J`b,
�:���D-����dK2|O����'p�H�`��O��$�O���'��S�`�<�㒓=�|x�K+B���G���<��O��d�O���P�L46�5?��5����G D�K<�I�J�0����g
/�?��)�Ī<I��E�:��� 	�(�L-㶄�4�Oh�'��'�r�?�y�([�f�V�C�N�cRp��u�<1,Op��O��]���>���d�9d>1�Z	R�X��?J>D��Fay"�O�4�	y��'Ny�O�)�vHKTK�;�t(���'�B�'���'��O��	��?a �Eg��T�^�{1R�����T��ݟ���b������O�KSl�������`�yn
��QJ�O2����7I�7m ?���Ƚdf��Sc�D��Z�bͺ�,K��b�9�?�-O��O���O0���O4�'9z�c�jF�*蓀$����O����O��$&���O���f�g������]�2>(��G�O��D8�D'��)UN87���(��HP�x�vyh�\7l�(�U��OE+v	և�?�V�.���<�'�?�%���:�ڶ^-K r!��*̀�?1���?�����dE}}�' r�'n �@3�R$J��1k�6|;$�j��Ģ<���?�M>!�^2}�����i�	v��� X)�򄖧S& 1Q7���e��i>)j��'��5�.��)�+l	B�)���U����ʟ���ɟ�	w�O����2i^=���{M\x3s�#��"�>I���?����'��d^�n��� kB��H�M��	�'(�'�j�H#�if�i��I�V�?�Y��ڨ(�X�)&H%/�{CMS%�'�Iş��Iџ��I�����>:.ĈҖF2������"��'F듗?���?�J~Γ4M�@#WH�`�p�e�w,�/O ��OړO1�2|�蝅p�R�a#�\8}�y;���3:�7MTHy���LƜ������$Ŵk��(�s
�HkRx3VJ��-�D��O����O4���O�ʓ<��	�4�X ��ah���=נQV�럀��G������O���t��k���T�d��N{��d�/��6�;?iP��@��i4�㼃e
�2�=�j�>]�@���ߟ��ڟ$�	��`�Iٟ�E�T�ɯrp,\�C���87�;�$[�?��?��Q������l�	O̓j�>L�A��X_|$��(IF��$�$�Iџ��	J
H�n�T~������D˖j��cؑ� ):D"�1��Iu?�H>�)O8���O&���O��KW�z�ʤ!��=��ݚ�F�O��D�<)�Y�8�'B�?m��
Ƈb͘)�W��a��<	/O���Od�O�c�v��gܲr�(��m]��9FkG�-� oZ���蟖ha�'��'IjL`�b95>\)"%g�_z��A��'d��'b�'�OB�ɐ�?�b�� �%�'Wb؝�v��~�Z���O����OF⟀�'�b�[� � ��k���(b��'G�(���i`�	�ED:P�r؟@�'/s�pr��`��JE
��t�����wyB�'�2�'�"�'��?��3�%I�DU �	�	�%S}��'���'.��y��'-�DJ�g�k�G��H��(IRj��!r�'{�'��O�BS�i.�$�H`�z���Oc�}�'�I�dz�Ƽ�"�������D�O���3�L���V�L�`�ue]*���d�O����OX�g���Wy2�'�<9���,�0=�7�B;C���1���<����?�K>ٗ	)j��q�V��H�  [bm��Z*k�x��K��(	�i>u�`�'[�ΓZ���E�<bۼ��7/dFjX�	韤��˟l�Is�O��dY{���w��2h*m����@f2,�>y)O��8���<�Qo�9Yk���΍�i�7i�֟��	ɟ@�əCx%m�g~aF�Q�]�'Wn���W�,d�~� e9Gph�I>	(Or�D�O����OF���O��p�*D46Ȫиa�5��͍cyb��>A���?i����<a��B�V��ܘ�h��4����d�O���.���!�|q���F�D%��� Q5��T�i�h��'� ����a?�I>y+Ol �D�@�1�����"�?"6�+p��O<���OD��Ox�ī<y]���IW�? lj6g�s�J�pPV04�,rD�'U���<������*�$ԳT�ݪ�1�e��>ix��x�i��Ɂ?̤�V�O�,�%?=λm�⍹�	�[򖌱gB�����؟��	̟���ɟ���j�O�xt�n��H�ɢ�-p�� ����?A�������	ʟ��<�T*@0^��j��B����a�K�|�I��T�i-7���R7M/?��¬��R�I�(�Ǜ�l�f�""G��?�D	!���<I��?A���?i�o��M�8p 	b�NZ�M�3�?	�����|}"�'u��'!�1?���G�ξW��glB�.����d�O��(��~z���0����T��|�FYȷ-K�UJ��7�H��z���O
�I>q�M�h�2|����	j�8�
��?����?����?yM~�)O����2N�(�u��-�($�fA�%M]���Ol�D�O��|�'M�N� �DȘ� ӂf���.ɘF�2�'��a��i���(&���i��HA,0�SK��m� ��'�8P�T���I�����՟��I쟌�υY��@�+#CM�JA0� @��w���ٟ\�����&?Y�I�Γ^�fH1S+\x�ʐ�ɓ8����ğT%�&?y�����y�����E��RR�����4!D~���^ʼ�)��O��O���|�����}��F�>{YpU�#m_�Bz7�'��':\���O|�d�O��V�|`^��7m+Li"[@nV�kE��x�'����%��kIץ)0���Q�EjZ˓]���Xp�Ѷ(M~"P	�O`�' 0��n�',�8��eX:C�����?���?���h��	�` ���̟pn�%�I�1� �dq}2�'M�'5�O:牒����!��Ap�mR�A�g6�D�O���O$�� p�Z�Ӻ���^��� L�?> ��A�8$>����Y�cT�O4��?���?1���?A�I^r�@Ab�y�.��J�`�(e*O~��'�r�'%��T�'x� ��e��d�g�4�����Q�������&�b>�����W���'��!� �j �[�v��s�]~yB�o����ɺw��'��I<;�x��g�J�+0�Pr�NG�n���	˟���H�	��ܕ'�@��?���܎	��ai��O��)�s$�7�?����'��������<�¨:5���F���tE �B���秊�'O��$\azJ~��w,j�
X�<�и�����Q���?����?����?A���*��$���f��;�bּ���1�'T��'e:�����O�b�8�d��� �q2�[�LV�T�q�=��O����O�,	�E|�N�s�^YQ�(�m��E��!�/+#d��v�H�j����X����4�����O�����f���Mϱq�Ȼp��9�R���O��t|�	jy�'��Ӕ)ߎ-�
���%��.vJʓ����O���8��~���#��ЁO���E����> X2�A̦;*O,����~�|"IH(~�LH P�DZP�I)��	M��'F"�'Y��4T�L`��|aj!�Ѧԛ5<n�(@�@:8��������Ɵ��?�)Ob�dQ�0�Yȳ�>�N�cc��8lH�d�O���	g���A��˓��� pص�5�T���O_TD�c$�'~� ��䟨���x�	Y�4k �	��OF#y�V\�Gc�g��I������&?�����ΓF6�)"�A��D�!�Ϲk�z��I���%��%?��f��A��\��DKR3{H�����hk<D�	9N�$a���'5��&�d�'���'���Rc�s"��C���)�$�'�'��Z� ��O^�$�O��D�Ck�l�t�μyXTa���qHr⟈�';B�'��'{rԸ�*�>}��D
�KF�[�K�X�l��+H'&�L�lI~�O�����y���bR���e�>D�p�k ˉ��?A��?)���?��Iq�\�$�F:1�(I�K�\��D��O��'[R�'���$}���i]\��P0�(8 �U�Ba�OV���O>���	6�??� ��~��	~�Q�jY">]m�HÚ#�� ���'��<����?	��?���?4�A�=�~$���Z�
�ͩ�O�?��Ve}Q����~�'+��1��''��S@��1wEJ�#*O�D�OؓO1���*�e�8)�lQ�4�� ����Ri B��6m�oyoΆJ� ������Ė��&e9�eP�yj��36/��H�R�d�Or���O�d�O˓��IΟ Z'E�>/?�HR�B�FG8J�W��h�	I����$�OF��`���4Txx��a�eB0θz��؉Tu7�"?)��h=<�I?�S���GB�X�ĠU�L�]�`Q`�@�	ş���ɟ�I͟XD�dB/}eh��.�<C\47`L�?���?&W�P�������r���l�� H�lQ�D V[;�&���I�����{��n�M~Zwˎ<�CH�af���(7���3���6�fVk�	Yy��'�B�'⫏�s�"Nu	`jN��@U���'h�U��r�O��$�OZ�<Z�-��)�F�`aM��fҮ�z�yy"Q�@�	Q�S�	�qf�4:ω�@6� S� yg�Y�֜� �T����f"�LP�	�9�m�⌌'������^4�%�I⟈��ٟ`�Iv�MyB��O� �k�LMW��:����Ym,�g�'��'�����<1�4�I��ċyh,B��̙������?1K\��MS�O`��b��zK|2�
�O?�	����Z���OKɟ��'_��'
��'B��'��ӣ5�z�z���F�,�vE\"O����'�2�'�R���'�23O��G�ÿ*$����ԓ7�\�s��'�b�|���D
*��6�O|�TG���Y��aQ<"j�պ��'wt���P��#2�|�Z���I`��6�@��K�e�����I̟���|y�G�>����?a��YR���E�(`$��`�B���}���P���I̟X$�\ʳH��vK�����V=�{r�wyۼ[��	׾iZ�i>Y��O��ɼHd�t��b��&�O�M��D�O���O���0ڧ�y�͖r!0���钐- �p3���?Y�P�d��۟(�Ij���y�nO$t�����nC�X������?A��?���z2��P�4����?
�RxI���u�hw��c�
&�n%/A�o��p$��'�'eB�'��'������,6L�p�M�*Д��P�HA�OR�D�O ��"�i�Ob�I� &ws�9�(T�w�6�Q��<A���?�H>�|B��؈Qɐ5̳iZA0��]6�l`��Lx~r胶(b&��	2pC�'c剐r�ܲd*cQn�h CHڥ��蟠�	ǟ��IX�'QF��yr.��<�ЄӇ�#�I+����?����'r�	џ��I�<iR��:,�� ���:Ppu�rF�=BZo�M~�%Ke���E��;��A���j��-�7LW�+O��iE�'���'�r�'�r�'�>����"� �__�a�w��(��I�`��Op���O�D"��="�t����P�P�QQ�+@�:�O���O>�ŵB^@7�5?�;"ʬP�L�	��u�P� 5� V�\��?ɰ+<�ļ<���?Y���?���i"�k��D���k���?A�����M}�\���	j�t���>���S�1d�4��\��<��������܄�0��6=?�MQ�hϡ2�LA�X�* %I�)����?�� �'z��'��`�I�!�fqKrl�+P�l��U�Z��\�I���Iϟ�&?��'�D��}m�c�%� �@���S��y��'[��'�O�˓�?I��mP*�q#���y#�A�2����?���kθD�޴����!蟬A�ʟ�Ћ3�[	!�B\��#�|h:ucC�'��ϟX����l���� ��H�Ԍʇ �B������G�o��IП��I֟l&?��	ޟHΓM����C`Y���m�� /�,0�I쟄&�0&?����ܦ���!�r��.�u�ѩ��Q�p�	9\��y؝Z �|%��i݁�'�?���M}�t�T��4S 8cJ״�?����?!��?���OS���'eb�'��m�c+ �b%�p�>�PFJ�r��':6mK�g`�d�O���G}�4��I�B(,)�T�Aq���@���F�'�rK����c������:��{�*�ə$�r5x�ÂnN�H��6)����O��$�O���:�'�y���,(��V"~2�駪4�?	�Z���	��0��Q���yr�\�wU���!k��_ؘ��&Ƈ6�?y���?���|x�D��4����,�[&���;T��/R<x*����df���f��������O��d�O����O��� _�>�J6	�;@~-k�oZ�4,B˓~<�	�������&?�,l�R�	%'T8dZĢ�H1>)�1�'A�'�ɧ�O�j����.-�d��t�؛>V��3�:�ź�O~�h��W"�?�uc6���<�uS>�
�3�Q�i�Z$�q�-�?Y���?)��?������w}��'h�h��"H�q#�4'za�0�'L��$�<���$�;( #�ꑗ5�LH"եڇ7�՘��i��	�j)�ț��O�ȁ&?�ϻ@H���+�#x�����.z�4����\������	��	T�O�(yB�)h\��&�)� � ��?���YC��XyR�'�1O����C�.��h��o��@ו|��'KR�'�t	H�i�	@=���5[J��.Y�[I �2�Q+�$>��<ͧ�?����?��*9x�:E�HJi���G)�?a����\}��'��'2�ә%�3cA��E;P 颎ĹQ2ʓ���O���O2H,2E�ȩ9��Y �)Q2	Q
	0 C�"8Y�y*���������lA��}{B�O�c�Oм{J 1	���HP����OD�$�Or���O<��2ʓ)����~�@��iá�dݩp���?���?����'�I�������K��
��u���S�d�Ɵ��I�_wZ�mZD~B��� h�a�9Ɣ[���2P��ڄ�^/���D�<Q���?)���?����?q͟ Y2f ��j���r�@�;=��e�ʷ>I���?����<)���yR	6W�	�aJO-u���c���?a������'xΕiڴ�~2�zj��v'�'kڨ�bC��?��`(hv��IW�Ity�O��k56�%X�,,���c1'�X�"�'��'8�ɇ��D�O|���O�$aeC��M��b�
���6�	Jy"�'n�|"�Ӭxn������YW�* cмR�	�SAd�Z���¦!���J�v?��'8L�W�]0|���2j,��h��?���?q��h�b�)� �`�$��H��=���OP�4X��'͜��?���?y�<Ox$��ʅ'<��p;�U���@��'m��'h�iK2��&���A�ᄺ;�4���q�m�*�V���E�>od��|�U���I��P�I؟��	��ː�+�p�Yq�\�K�V�ayң�>1��?a����?iP/�n���A�&|���ߗ��D�O��+��I�$ElN�Pt%�Fx���`IA �����@:�	� h�y��'�t@&�|�'��P:u�?KD�#�JW+Yg2h�S�'���'�"�'��Y�l��O�$�Cir���T�G�P\��j����OX�Ȗ'hB�'���'�V|�U�R�!���U�[�z^N�#@�i��	�o+�=�C����jۮF�a���O�eh*ɔ������֟��I��<�I���D�o�b?�0�G�-ĭ� ���?��?��S�$�I�\��E�`޵��+��^���E�A��" '���IƟ0�	�[<l�a~���w��u��GZ,W#l8�ߛ��$�k֟�r%�|R[���쟔�	�� )�fH���ռ�
%d�ߟ��	vyB�>��?�������J�A1�Wq� �Ʀ
`u�_y��'��|J?��Bŝ( �&uY�f�<?Qx�0�IT�DВ�U�p���z2��O��J>a��*�Ĭ;'-��uaT��sM�?a���?����?aM~R-O���I�0��s�k� j=�Q�H�-����OD���O:�$�'�b��nn�)�CIѹ> ���F�F�IF�|lZd~�f/:���S ~���5�h�J��S�O�^@�
���(��<q��?����?���?A͟x�HG��8�8)��CDϒ93K�>q���?!��䧝?��y�a�(,�PS�̞�!�j���?��������6�Oȑ�5��t���� ,Mb�'P��ӑ�m�6� �����O*����Px��b�&9ǈ����<���O����O��,��DyR�'���a�F��);�bF�: ����<���?yI>�*�|��;T�!49��{�[���P���x(t�];i����p�l��IEB������k%�@�O�M���$�O��D�O���$�'�y�ڹop��`T���1��]+�E���?��U���	ٟh��d���y"d�0m
M�4(bb �ȫ�?	���?���=�F�ش��Ċ�0 ��)���uا G�,#��N!.���87�����$�O:��O��d�OZ���9Hp��+���`���Ȝ'�6�!�I��d�����%?牽G�^5)��V��-s�C
3
�4��'6��'�ɧ�Od��	��Ѿi��+v�V�e���3gC.:��OTu�fN[��?�-�$�<I��Ŏe| ̱�Ŝt�:`�ch#�?1��?���?)������i}2O|�FfR#�=��I$q4Pyq'�'BR��<����$@���:���!���Qa*1U����i��	���,��O�M$?	λk�V��Æ9C�D���)\$����ܟ��I͟���ϟ��Im�OB��q)O�RZpe­~�|r(O\��H^}��'8��'F1O�ɡ��
�B��ŋ\>Y�4�`��|��'s�IoLou~�@:�D�+B%t�.48�E�o҅9�,՟@B��|�\���	ٟ��	���3D#Q�K0ܝ�0N�bV�]a��G���Imy�A�>�)O���*��͝�`@�!�q%TAϺ�@��cyRR����ӟx$��O����CY�j`��Aa�3Q �c�K�&�F �fD~��OZ\��I0)�'Y�i�HaJ�ꑀE�(b�B&�'b�'!r�'��O�	:�?��h��B����0ꂬ����c��㟸�I�P��|������ODEA�+w2����2C�
��m�<�T!��M+�O$
sg�.���!��	���<�C��4@Cֽ�"P۟�'�r�'M�'���'��S��hC�Ƒp����	�	<��}�'6��'�����'�;O��;W�܉`5����	��q��'U�|���d��4���O�4���m	��:��!����1�'ɼ ن�[�8BA�|�Q��S�d*��6rm���3o��hb���ߟ������syR�>A���?���x��E�����R`x�$Z�1�����T�D�I��&�DJ#i3Z�ұ�2Ie~�1��DByBKG4j�(� �Ø%�O�,��	%��$N܊�1��!K��a��%�c���'��'��S�<Q� T����f�����t�&g���$�Ob���O��0���<��+�1u,bX"�ˉ  ���������ş(�I��r o_~�-(�����+�-�
 K�tcqō)��p��LRe�	iyB�'g��'���'��'q�L��V����h��Ʌ����OX���O�������b}�
õH�VСe.��;����?Y����Ş�4��G%�|Xl-) ȁ
�|�����M�_�P��G��8��$?��<�*
cID]����&� ]��9�?!��?��?�����	m}�'�4a�Un��z�+4��$� ����'�b�$�<���?a�'��X��R:Ix�X&�D1Z�U����M#�O�h�U�J9�����d4�x�3͗�,T:6�,�����'��'�B�' r�'�>� ��U��%Lg�yчw�n��_���	?���Oh�D�O�c��cN�&^��D�T�X�W[�hz�j"���OH���OVx�	bӐ�
�d�3�o����9A�K^�*x�+�&��S���������4����O�� �̈��n�N-z0yC��)ef���O��M�Iӟ��I̟��O-�Y��N� �
���!4��!�.Ob��?����S���8�8Y�7��%bd�ag�;V�L��A>y-��3�O��	B��?�gb,�d�� 8��rB��m��q�mC�8�����O��d�O���)��< �'�8� �Aκ8aL91�����?���?��^�t���uN���C  |�	�c&F�n]|��'s�Aa԰i\�	:
�(��Ocb��O� \1�����c�E�/f�U	�����O����O
�$�OZ�,�#,\�[^���G.Y�E�ܜ�&&��$�O��D�O��?)�I�<I���)!����=6�!T�����{��r��L�anZn?�eo)Mо}!%�G\�0�e	 ԟ�Ҥ�[SWbLq��RyB�'��Ȁ|A�eA�+N�EP�E�͞}!B�'�b�'�I���d�O0���O��t����6lˆ\���5� �	wyb�'���|b�Z�qE�����9U�<� ���5U��	3�T��B̚��L~���h�<%���ɴE[*5!a#"�l���؟���۟��Il�O��D �SN�8�/�([C��G'׎ie��>	���?!����'i�dZX}J<Z�DM��*��K���'���'�� �4�i���z�J�!�O뎚�|m�Y�bOՕq<�;B��'�'��ğ����4�Iٟ�	�$�(�l��Pǆ�k�(ߞU�8�'듼?A��?�J~J����i3i^)L�$�89D-�/O���O�O1�b���eX�U�&T�J��؆ŏ2.�V��H��?3���s�Zy��9C���E��*i�A�BF�2�'}b�'M��'�����D�OiI����P���@���:}6T@0��O��:�IXy��'�2?O�*��;B~�� �7	����6@����,`4��
3��d��g��ì��tYRu���A�!��O(�D�O���O"���O�#|J7��r�L8�������a��\�	Ɵ���O��'�?	�y���f;t�3"m׷(��8I�� ���?I/O�
ujb�d�la�y;����VK�4��*R.Cbx��_
5����N#����d�OF�d�O���ӊd?|�o�vҰ���i���d�O@ʓ\�I柌�Iٟ�O,���?��4���Q�WHdA*O6ʓ�?A���S�)��H�@���{(�0�3ea"y�D��n`U��O��)��?��I ���j�c���EnMy�@�!��$�O���OL�d5���<1G�'��cS�D�"ľ(qW�:H�������O"㟔�'�� /�, �׹c˒��Pf�";�b�'n���Źiq��9%�Ƌ<��
�0ţDi�Ā9��e�%��d�<	��?���?Y��?�ɟ�I�����sĦ��AػZ�$R���>���?����䧌?����yRHL('��}�t��w��H�/��?q������ڤN뛦�O�i2(ݵaj8����D�����'�҅6ƃퟴK�|V�|�	���ؿU1����ް�B�%L۟����p��ayҪ�>����?1��qX�$��1Gf�d�g+Q1+�� ���W�h��S�-V  id(=3���3	C�� �A+O�l����BʀT��,�)�&�?��!m��#�π�7�|!ri��R�R�z��OF���O��$�OТ}b�'�X(�#P'yF�1'�L��k�������I۟ �?�'"`<�G1:�I�w��	�LE���?����?��D�)�M�O����B�I�3vn����@�Hph� S'�x��K>I/O��$�Ox���Ol���O���U��,$�mɁ�o�a�B�<�TW����ڟ �Iu��4S~%$���>%�	F�I�k�`Q�+Oz�$�O��O1��� b�7l$�M�<�d���2n��`)㗟��a!�0e����M��qyb�Wr�A�#�gm�W��'���'��'B�����O�`Bd�ȥV��$��(Ġz]
I�w��O��-��Ry�'�?O�dҀ�^B��Δ�SMȭ�3	�
%���<!�N�"����@�S��[��@�g�B1:���U�~��������I�4�	�\�I��F��ݍ$���w �q�b��tb��?q���?i^�|��ӟ@��k̓[T�b�*_[:��0�x��&����ߟ��I�Gp�o\~��m�$�'I�<z"�K5��x�k1@ӟ�C��|]��S�l���pc�Q�8F���`�%������I}y�>��?�����i�0%j�ه��s���as.ؘU��Ieyr�'^�O�'�e
5J2�U��O�j�-����J�нCrGP5h��ʓ�׮�O�E�K>G��,�VhpcC�Cx)Hd$���?a��?����?�K~+Oz��ɠ] >}WZ)f:)�|�$�<Y����'��ן��s�ِ���Qp!�����"Ee�ş,�I(~@*�lo~�d�nkP�~
��:H�bA�PDg����&
����'X"�'���'���'��3� r�3�%�82_tqbvk�'��ً��>���?	���'�?���y��,��%�B�b���Y�]4�?������'7��X�4�~↗�_�x׫V�] $�p�l�?���~�b��i��~yb�'&�eZ-q�0L{��Ɩ>��(u�\"s.r�'"b�'�"����O��D�O����$��z��Eo��r���¤(�	Uy�'��|��,x�j�)]4o1Pd1A��|��ɧt��)Ф�G�wM*��|����O�T��'��i{�̆T-Tx��G���Tq���?I��?)��h���ɚUT��Y1&ܑx�̂2
3V���CS}W�$��F��yB���X��ᛆF/��Y���?����?���sX��ڴ���J#w�ؤY����k�OQ>�L3�dQ<J���|�T���I����	֟��	͟ Pc�=o�Ҧ�B�4�8r�*�ny�>Q��?�����?�F�F� MB k����ũ��_����O��2��I]M��X�ÔU�F�&��dMrQV�%[T\˓{�&5qq��OxQ9M>i)OL�j Ê�	2�X��͙��x�Ä�Ox���O��d�OZ�$�<qX���	H�n� �j1�`&��D��ɟ��?Y(O�5?Q��p�b�K�)��cq�OZ�Xl�Y~r�E8?qB���:T�O�#s������ƩF膤��*F3"P��'w��'�B�'���S}"�p`A�/s,���m�/
����O��S}"T����v�xBJ}Aᇿd(ԕ���q%�$�����$�	;O�ln�a~� ��RP$�hvaP���ͳ�&%�&�r�n�̟L�Q�|�^�b>�I�s�LL� ��]�=+!/X
h�0��OD��O��9��%��E�Q���a),� �TBy�[��I�0���Oâ@d�֟z���̑�'֬�6l�>Jm���Ϋ�����B���?�`�OHȡ�o�V(&Az�c��5���O>�$�O��D�O.��P�-\r.E��HP�R:)\ă䮙��?q���?9����?�+O��ĝ����	<��2c�� /�2���O�({C!a���Ӻc􉞔�bc�1ʃ���a��vΜ�h��9��F���ȕ'/r�'���'�b�'��ӏ8:=�s�B"N;hpu)��jD�'r�'$����'7�7Oh��B�ȫ=$�	�o:�J��D�'D�|B�����2כ&�O�ewG�A}xq�F8J�^=��'u�Y�A֟���|�V�D��ܟ��r+�F���N�#�6�S�k�͟L�I��x��my�e�>����?��
�X1A炠 оTA���Eh�K>����O�$$�� ���S�B��ۆ"R�g��ʓ �}��h��M+���T��?1�'���& λ%u�!�p	$fB@U����?���?���h��I%�t�{!-�	��B��P[���O�(�'���'wr�|R�'i�M�ih��C��5=n�[D� :T��'���'1�K�i��iݡZ���?͙��;a�� � ӣiz�xB�Ϡc0�'�I̟��Iӟ�������I�� d��@ΊQI� @<~K�x�'I^��?���?aH~���C�N)���͠\/P �stz��/Or�$�OʓO1��tbRǆT%(�X�䍌Pil�qS��52 (���<��F�o���������"`X����%�� C�vF��$�Of�D�O����O<ʓ��Iԟt�UI�~��!��ڙ7�P�j  Iҟ��	P�П��'��'@��B�����
+@�a��I�|�ði���$$eS$�Oir�'?%�;?4�R)��T�А��� ��H���d��؟��	���^�O���i��/����2�0@\�����?���
��������ܟD�<��+ @�@@�����5�Lq�6��T�ʟ���֟����B���'Zd)��@s-.�Pj�/>�1f�J$C�0����'G�i>��I͟����6@�i��� DG}(��Do$��Iݟx�'t���?����?�ɟ�� �'L��w�:#���S���'c��'ɧ�$;�pJ%�͒d;)�j�+OJ@bMQ6"�,f����S l@�̊C�I���`�T@R�RV�����^8D�	ß��	֟��	H�ByҦ�Oy�%M�Wl�t �#��U)�'���'&��d�<	��H�j�І$_Ȥ0H�'��jW����?�!��M��O�!i 'v��D�S�7����@�:y~P��ӸM�F�d�<����?���?����?qΟ�[�#t���[�H��I�<}�j�>���?�����<����y2�[ƒl� ��;����s!L�?�������'7}h,q�4�~Ҡ�IȘ��_��t��o�?I��	d}8��O����4�����?F��L�U�D�1�HY�5&ʣ-$h�D�O����Oʓ�����	�DI�.܊9��(�GСIRU����l���d�O���1�d�<|�,�7p ��ru+$'�˓ܨ�F��7D0�(���� Q=OhU)��=&ޤ�,D��0�'b�'�b�'�>e͓o`�����|i�G �*E����$�O����O��hΓc]��:�j�ԅ�(M
���s(U������	� �z�o�n~�J	2u��O��y�� �dD9�� ��9O�1#K>�,O��D�O>��OJ���OJ� �]G�"F��iY �Վqab�T���O���O>�$7�)�OrtHHISx
�%�ύL6�d:6��<)��?�J>�|�$��z2тQ��
Q*�zŕ;l",kٴ���@�|���'1�'?�	�S�6l��F��(M�2��!v�`�	�������	ܟ̗'��ꓹy�%�1J��_�l"�.��?����'�����I�<93���־�JDC(������$o��n�L~r*�>�@E�0�r�
�n�oN�� B�C�o��aٲ�'�r�'���'B"�'>����k�⑐G��- �4��U
�O����O�d�'���'���OI{ � �>2�v��ց�#��'���'��'�u������Io��
R� �v�n���H�"Z��en�/!q pR��G	}�>�U8X򾭲҆ {�T�p�j�K!�Q#�l�%5Yإ+�Q2Rİ��3W�E��M�kΚ��JU.��҆
\/Y}��&-
�eZ�d�%��%{��%2�H��\z��Y$}�����(�3=2�h����;sOn��-�5w� ��Х�����7e��K�*�v�T�i�ȪP��1ggęSe�T1IW�����N�[^6�p�ʒ$o��r��Ǧa�6��&�=�9�Y+}?"�z�E�wf0Rȗ.{:�����B1	�15Ԝ�z^<�q3r
I�x�(��`�xM�2)��
�XT"	�g�9K*���#ꉓA��T��Dհ>����� @�f���N����㇝�S�L�,%(��DO�g��X�Ԗz_�0`�	I5A�����Fɏ2 `)9��	|��$����x�LH��ix� 6L?U��8@A&�.��ge�*@��;F��R:�D��j��B"�a���i�0��eL���J�`��Y{Ǐ�F��@@I�,y7��U&"L�1 ��9�ď1BA���D9|�&h����O����O@	�'@���pAT$��e�G� �69H��'��'���'Y�'��(U��Y@4͕�|����� @���1�Jޟ��I�M[��?���?)7Z���'���V��NYH����5t�e��'��$��'_�'&�S)e�*����ibҐ'﶐06CO��֠I�I
�M���?a��?	�\���'i"<Oʬqui\����&AY�<vt��K�0��o��D�O����O,E�%�l`"�5��@��OR���O^<�'��͟0$��r��B�mt΁8�n�	qg�D�s)�Qy��Q�>$�b�y��'���'��S)o�D=� ���%p$��1'ԻG�T�DC}rQ���IR�	蟨�	nkD��(H72ז����p� � �DP���؄�v�p����0�	w�S��MG��"�	���H���ȟ4�')�|r�'(b��:["��('�萋�.ϐW9@��U�r��}��'��'�r��m�~�j*��jT��3|Jf�Idc߬1����?�N>����?�	\Ř'�b�kQɔ�nM������(|�;��?���@�Beϓ�?)fY?�	ԟ��I�nչ���"
��!Ǌ��'����ʟ H�N�\���t
�����YF, |�1j��*�?IFa�<��I��f�'���'��ſ>A��[:8�t��uJD�oO|��	��?����?�$�o�'��!,���L������קs��XP�N�ϟ���Ms��?���?QtS�\�'E"q��a_��������M��'��@r��d�|2n�<	�#��i�׆%�Ҝ��m۔B6��Ըi]��'rR�'V����O��I9$l 9�*J�(����`nM�N��⟜�A؟$���j���Iӟ��\e,��,%d�a;F�:8�L������	��S�4�|bK�T��y�� ��60r4�+(�' r(ɔ�y��'"B�'y��?�I!������K1�d��FT�	ן���M�IWyR��a��u�ݡ{��)Z6��#f���'5 �A�O��'�B,O��SCp6��5�	$�x����[ws��$�O���/�Iҟ�'&t�y`
S��%�u/ʪFV4�[�e�\��Ob�d�O����<(����1v�T�QA��!��!QD��&(��d=������'7n�YL� S�"J�4��"Ōg��İc��O��O�1��<�-�����O��݉?{t)P�"X�YzF b'��9WJ�OD��<)R��t�'�����)֢<������Д0�`Ѫ5�'a��1D_���I������d�Iy�̜y�fŢTޙi�t�8�
>3"�'���U�#<�'f�1��F	���ђȍ�_"��͗����O
�D�O0���O,�S���xD�K]�kZҬB��F�	o剓
*P"<ͧR���͓�?�����(?d|�s�E4�Θ�'��YI�6�'r��'��E)�?e͓1L�x�g�O�&kX O�t��̟�$���I�i ��?��w�*pZ��;lܔ��MI45~u����?�����|ډ�bӌ~JdIk��4>@A���#�'���@���y��'��'J��l(����9�F��)Df��[B��ϟ��Iw�Oy�-
f7�%�V�E��Ic� P���'w�)�O��$�O�i�<�O�b�JB�����e�+;L�����?)���'r]�,*�L��!"���
5СI$ ��3J���Mu���I˟���V� ��I�O�у��o�nUaD�Ŷ���jD��O ��6���<�'�?�ʟ�ꚨqR\�!��fv��D�'�2�'��-��'E��~���?)�w����PJ�<ݮ%�v*׹D�:$S)O��Ļ<I���?�J~Γ#T��e��}���pG N�y�(��/�X���?������'���'��T8�x�Y�d�%�۾+��æ�O���?����'��Iޕc��� ���DHAf�����,��8�`H��'�rg|�>���O����O>�'����@��y�G퓻D��ұ�ܶe2����Ob��OʓO�I��b���O����\�c����oPD[�����A�������\�Oʓ�?!�'Մ�J��,J<xDpv��D�~�A+O*�e����K^t4ͧ�?���?A�C �VU�נ9y���熠�?	���?Q�Y���'��Q��̻yع`v�
/�"�8��'j�D��'[`��'bV���'��'���y��I*t4�䂅)^� �k#hĪLW�>a(Ol��<i���?���-ެ9#��V3	I�͂ᕷF*(�A,�<Qg�<���?����n��T(����(�t�^\T� �gi�?�)O���<���?��~�<���}�0'Â[���C�$�g#������?q��?����(�@$�O,�Δ���ɻeLց���g,U�[��'�����I� ��h`��O�� �gb�'0�d��Z�҅��'��'��1Z�'���~��?I�T E+S���7^����g�rTQ/O|�d�O��Н%��D�OB˓��DOF�e�b��
ץ����ׯ�?���<���&�'=b�'Vb-�>�!�E�'�y�ޢ�5�p���?1���?I�g��<aO>�)�(4����H���j�.�j �UK�>t�D�O�]m�ǟD��Ο�����D�<Yr��6^zAz�*_�>�P$c�N��?1�˂s~�Z���O��\��O"҉��8���3GH���U7��6��O6�D�O"�$ Q}2Q�����<Ib��$m�b�G*I 
�+֨��L�	ay�Ȍ��yҦ�����'�=��9K5��L�^1����/|�`�W�'���'�����D�O4��y��6Z��E�$?G��9��Ҏ�?��?4hΓH��ϓ�?I��?y+� �3v���(O�q�G�-b����O(��'�����'�R�'�R�L�q"9�"Ċ$f����	Ñ��	�'�R�9�'���'8r��� ��B�{N ��1`T7`�Q�',�؟��'-��'cҁ��y�"I�v,���Ț1�dZ��G��l9���'�"�'!B�O.哅����O^�)�(\�gJ���Ǜ0T�dtH�(�O �Ķ<���?	�`)28�'�$���}�QD�)26r�b�S�d1��'r��ؖ�y��'H��'�?���?����$���S�Qm�)r�d�����OD���O:�11����'���I�*p6�P�hK0�<�@T�)Li�ܷ�y��'s�6��O���O��dT}�ș�$�6�4%��#s�
(@�FB��'Rb�Y=�O�ʧ^12�Z�
ҪQp�����2P{�#߼�?1���V�'n"�'��/5�ɩM�̑`P�1G�������ɠd����	o�II�D�]��y�'1r<��.�y������2&���DCg�z�$�Ox���O���>9���yR≋�t��#�΋nnx���ͻ�?1I>�pd�<і���<����?����@��
k��i��[�Y�QC��?���j�'�r�'��'�(���&W��l���@�>e�|!pS�<s�f�0	r���������l�t H�q4&I�AG�{�)���?�p���O�O����O�T�ǈϮMJڼ"�
:l=NXQLA�=���MV�D�O���Oܒ������9=ą!��A#�Z��C�4�ؓO��d"���O��Ӫ�������<��l8nb�9u�R Z��} �2O��d�O~��&�)K[�T�'x��ۇ'ڑ?]��r抏X���j0�'|"�'R�I�Q�����v�G�	��H��˳-b�ͱ�H�O\��OB� �9O^���H��'���',H�86�L�4��f�@�6<td�0�|r�'=b�~�"�|"1�j8��\�1t��R�$�5^P,��'U0��'J�ne�Z���O��D�O*��'��B�R��Ȼ+V�}P�����?��Z>H|������IX:VO���PB��7ٚ�r�mޏS�&x����Ox�$�����ğ�	ןĩM<1����Y�1ò�c�����
�O��H�%�O��O�˧!�1��?ه����t�2��4L|��d٨���'^��'��1�$�O:�Dy�4���F�6�d�Hr�K�4�����Ob�O.��r5O����5O��D�O���3)��i�m->Y�Q)"�$���O��P�����}�0{�pĊdD�2���Je(�8h�'�L(��'��[�'���'���?�S5+@"jx T�.�e�D�!��O�)&�(��՟�'�,��՟\��`
��z���n�ujᣚ]�,��8n�	ꟸ�	�� &?Y���E%Dpt��AI��,
8��<���hO>ʓ�?�R,NrtG!�8����!=:�Γ�?����?!L~��[?1�I9/X4A%4_�dYQB�G�_!��	˟�'r�'-�`���y��'e��T�܌$�W����ǀer�'B���y��'4�ꧯ?i���?aḟc�x�8��P�o�	�2�L5����Ot�D�Od-�є��'M�S?`���vk�=��h0��ɦp7�I֡�y��'I�6��O*���O��$�S}�i^1/��3V�d�@��i@�4��'�^����<),��1����DY3�ؓ&cp��4HN�A�b�d�O0mZ���	̟��ɾ��D�<��(��#��e#g�ς6��#�JW/�?i7��<QK>!*�$]��3O���Z�����kp�J6���l��p�	����	����<����y2�G4|�0��I�(*&Z��H�?q����DǴ]���`��	�O,�$�O�� N�;Eˇ���:��-`����'���'x.듰��O���y��]�kd�1��c-�d-8@-B���!]\��
wf����O��$�O�9O�5)� ?�$�*5��+���"�O��'��	���'�2�'�R�F).����&��)q��x0%bE�J�T<�'E�d�P�'G�'��[>�	�ܓ��0cC��C�ꆹZ�R9�v���$������g����'H���샎0F��u�\�i}N4B�+��kz�S�'B�'�B��T��~*�R%2�U,g�d��C�ƕ(�$�����?�N>����OdM��|�$Q��	��al�pc�'�2�'a����'��f�~���?i�H�6�8��PO�|��A�/��qN>��0=��['��� iEsWP��C��B��s� �	��M3���?���?a"W�XH`D;>P�2��t�4���OD�$�Oqy��Q�4$�"@�Y��M2Gr���pg�5W�����'�hx�`�d�O\���O� '���I-9 D���5G�^,S�n�1����ɥ2�#<�*�hT�@1O����1X ) �	�ZcT�����<�����O���?a/O�ʓ�?�'����T ��h]��4L٢0�|#�G`�'[�TF�=�yr�'N��'��pQŹG9t]�!��7AX�L�0�'!��'��OHʧ�?�*OJ�!���,��p�-�)t����"�<��h��<ՁP�<����?A���B�OV���g`J�!R�<�dA�6,\!P����d�O��d�O�O��Di�0��%��}���	�`��\s���c��O��!0Ć'_����O����O���^=�@�@y8S@�(�OG(&T��?���䓰?��#q.���gi~ų�O~�$pTh�r��a	h���IΟ|�	G�S�����O��Z��xtΙ�p@��>:�('��O���>���O����(`gqO��i'�9Ea�E3g�W*��$��'B�'x�X�'����~����?	�e��14�R�G��y��	�AД�H>����?���^���TbW�|���lQ�jRE��$�?9Γ�<���4H�v�'"�'�i�<�%=@�I�$ݚc�A��I�ğ��I۟t��5��򩝠W�aȄƀ��(��F0<�@�	�O����O����O&���On�����s�$٠HNs�zlatM_�r�^ʓF�2�Ex�O�H�A�'RC��0*
-"%����O�n��6m�OD�$�O~�d�Z�	I��'Z��Ȅ��3T�}r��#$E�(`�$D����Nx���O���Oy�!��h/��9�$_�`,����O����O�˓����O��O�y���Ap�Y��Õ�1n�:�.�$JN�H�Q���w�ˎ*t4Y�G�	�<�ءB�Ǫ,Ę�"��
,p�+D�#�X�:ҁN<\5v'a��?I��?�����&����!$C��:�{v��x?��P��M��y���'R�'�'��	`�,�#��>�85�p,�/1�@̠�H?\�t�A�V��
)�b��t�|!c�"�H�J�.�%%�l�GM7v��R�9ㆰƈKU�,!�n�.{ը̣��0w�Д�4H=b�^9��7��P�G�NA�|��Z�z�Ǩ�ar:82��G�X���ؗ,�k�����$�,YL��	�w�
9PF��uZj���L�t�(�*�_ET�R�"j,�*�%4a�j���� !/o��Baעhl�s�(�c}$@2(~^��5 ܣM�ؼ�%`AR��9�b*��H���:�E�yh�Q4��%��̟T��gy��'"R;�X�oR8c��їM)������z�m�4m�n��(wx�,�w#�Z�Rl�!�̦DY�T��g�|�24�H?��+#]Ax��*4�lӎ@Q �	.�tH�fG܄Yɦ ��؟4D{��	0 {�9���+�ƬQ���5��C�ɾa�FM�7�_�0��h޺.kz�'ABꓢ�Y�s{���'qr�i�  ��K�4Av�9��Z�DTVq#Eɣ<Q���?Y�P�0�!�@"�� ��\�R�Zw�@�7Sje��E�Df��(����:�8 ���
�ΐ{``�?A�2�װK(�Eq��@85����.�"����	��X$>1 hX�3�b1ϛ�]a y�k0}��'� ��$U ^GZ�[�H��Tg�X��P)�� 	�~��I��{F��� c^�na�'e�9`�k�>����䧨?�ܴo��
�]g�4I'���\���'p�Ѕ�ދd�@q�bv}*�f�8:Pa�9p��#�5}_��#P�����CV�vq�����0|2�/�Q?�5�2	:i��QW�\F}���?�������4S�dj��_�~��E97	˅[��A� #D����%�?M���r�˦�F��0�	Ш��u��-"5 �e��s����R�O(��O�����M��U����PyB�i��	Di�Pj0C�n�	rᔌCS������9O2�(
V�R�3�	�.�8����
�b�piÑn���q��>�-Y|u��ǒ��}®A0l8��j�vܞ��o��~�0︡�I�,D{��'�Y)U��h���j����wt��ȓs��@�H�|��P�R/�}�L��:ő��'��L3��T90��&��mc6�Z8^�xQWH��1������	kyr�'��8�&5J�iP@�EG;`�*\R!��U������xmڱ'��s���yK0t�ã�!���$A�cK�� �i�$ꁰ��x��*)���X�KDH<y&�d�֐AW%#��p�e%^q�<�WeΑy)�����'�b�`uL�b�$�`�=^��#�i���'�f�U%T &�x%�K�+�*�1���	8�~��?���?y%���?��yZw��RS�`:�pR��Z?*r����DX�t!�>ӳ�A3@���CN�Y�2�2�c �6	���[�P�, c���
C��<����'�R��ȓj/T��2�X��L�A�޲` �i���7�~bf��e�� ��n� C����X���	�Q�Sݴ�?�����?q۴3�tqЀ��;t�t4�wF��Xؑ:s�'ȸ:t�I;\	��O�Y�S	b���a�,1���W.�;5f�LqV�qo%��S�O�B3��6(	�QI�d�D����O�EIp�'���' ��S���p��Ϩ^+�(9č3K�:�'���'2��r!':oHXYf�߉[l��@��$�W�O������ u�V�АɑFl�0��OT���O~dڔ ������,��Ky�iY�I�g�2Oz����HM_Ɣ
O<i���H؞�3p�B�r'�=y���g�n4am:��=�a{B���zm�׬�u=B�P�ȋ��&�z��ISX���&+��M��
�e�U�P���6D�����??�y���O*q�7���l����X9���tH�9�jyX���4�f��g�K��M����?�������O��n>�J�y�LM� �ʅ�9\�����$�a�����M� >K�b���W[.����Ey؟���a�쉚V��)wd��@�Ô�M>N�cc��kH<I�jô ��g@׉,�8����v�<�g�S�o��8��� {b�"�
�v���X�[���b#�ip�'ߛV��0T+:=�Nܙsu���	��g�˓�?I��?�G�ؑ�?A�yZw���2h]�W��M�����4bl���d��w��>5�ץ!b�鶪ڦ��z�	:�-����v�~*N!h䋁�+�d8k�Μ�[w��ȓY��țS-ҷ[<
좑i�4������~"D�%R���\�Iʞ����,b T1޴�?����'�?�ߴC�҉H��A	���F� �I:4�'��H���'`1O�3�$Y�zVn�;'����
�a�aܲ"'�	�c>#<E�@]��~�c�^2DsPHd�����3�r��M��y�^�H��Q8��K4�B��,8���v�J!Zk�U��(]I��>y�SF0�E͛�p������ZX�C䉾\4ls�JQ�{t>Tr�ŝ�CӦC��9xlz���j���+sʡ�7FF�xf��IQ��O����q���C9xq�͜%*{D] P�;D��:�O�.D9�!�<r<�i�D9D���M�Rl�$�p�U�����7D�d c��,T�����*��DE��2A)D�@Rs�۩=�X@ ���z�tep�'D��e��.0VQ ��J*u�8��6D����݅]��(�&�"��J5D��+��C�|�f]��&��R�qu�3D��#�"OT�qt���D�ǃ0D�ðț�X��J4�Z$�T
@b/D�Xk6��P\0ʇ>p���!&1D�IF�K�_V�`�dÛ,A�V�+'C:D�l���
��4m���b�Q��;D���5�:e�:�w��Hv� �#D��4i�4��Ed��6�V<��'D�$�$�=�Q��,.�ĚE�%D��1+Gt�⡈��������a'D�Xr�"\,[�@ԀEcBW��pl$D� St�%��U����V�ɉ!�D�i�~��%IE=l�0����!�d	PzeR'��Is����E�O�!�$I�m],�KM,	o`�l�ݏFe!�$��&��}#�O��y���2sG�?�!�Z{��p����0��[�E�}h!��  X'm)
c�Xŋ�X��S "O<�YV득~,�)�����3"O�ɢ�&�ihv�8.�Zo&�h�*O���� D�VӼ\�A'N�<cj]�'�J�9�� )/�A*�'F	1C̩��'�T՛���hmR��$��<:*�b�'��	Q�#N$Q��ptL��8�(�'�`Qf�$����&��C]J
�'?����͙�4�q	v���8��'zLPp���*"�̛%O�)�:R�'��!O�� �őt��j�|Uz�'7nQx�c�RЙ;�� |� �z�'�j�P�(X�*�0���I��,$�R�'g@!(W�V�K"L�����9q$ҁ��'��9����#���G���;�8�`�'0$)�1ԁU��ZټL^��''��2W�'5'\�BՈ�:^U�5�'�����~��DO�(�@�ȓ_ʴ-�q�[�~���X��r^��ȓ`�X1�G��-=���I�
vo����4%�]�g��<9i�ݩw�Z�"����ȓjJ��d��w���rB�S}�d��U��m#����<�´��:�مȓi�ޱPƍ�,���2wE�v'H��5�yv�ǔ���G�ۉ�$��+���&�#!��s�*UPT���ȓ6j��t�3@�*u��'�W�m��3�)
c+F!t���gVQv�,�ȓ\[�	�G��9L�J��e�R�GU�<I�&�d]p��qC��K��<�6 �U�<ѲC�c\-�Vʘ:,���)�K�<���R�w�\���F�b49x�_�<I��ܤ�p(2�
������Y�<�$��#�r�����a.��t��T�<1R�"H��#�X�ZN�:�\�<����Ji�u#��G�2[$(c�dZ�<��f� �*��t����:`Xs�<�%�D{��!W�ĬIe�Ā��Ei�<�!�}V�<3�n�+`G�<����k�<Fg�'$"��w� &^�I��ٟdsR��qO?aׯ�
pS`�r�&.�8�z�E�S�<هK
���x��! ��*E��W?	�gY��v4LOF�B񤞄@�xZؔ�f�K��'a�E��ƻf�N�Z���\	���5�
+
j����S����ē�Ќ��f�%uOx�R��Ť7_���>y��b�(DjcJ��g��5��4�vD���ģ:eV�#a��y�k��DwT���S�?��d�$��i�,x��;4��-Ɵ����Y�<j��B�N��xq"�
%a��\���/lOP�L��۱3;��E��!$5^}��9��+��^�H<��#�$�� �'����tԉ,NL�`2𠈑�{��zU�ز�]��2a��l�iA���U�n��T�1����瀌,G�U��J�IG!�dš:��	9񎏚d���q��Вn�X ��-�?A�/�G.9�)#?��-y�Nϛe���a\SI�aλV�VrreO�P�b@%�
=J|����P�r!�W83�L�Ч�̤tΐдb�%k�v�K��~��t�'LO(�Q���W90�X��'J̥���]�Tk3��,V�=�`jؖM�,�kG�&�jo�`�� 
2eB%�r)�z����t��#ѯG�^���ς�n��1Q':�lԃA�u�<�,��5Eb	�&���;Ћ�),��h���!�y�.���l����K�S��(B�Tf��CT�WR�27&#M�"��$��'+*Mi@��8\ܨC�j��J�0�s
�/�Y����h��l���2QTR%�Ra��q��JM����2)�m�`�5j��Hx`
�RR\ϻk�ά����& �јf��j�^M���5P�2l��&$0ꔅI"`�yjh�k��W��E�N�'�h ��%�^bu��%4����`H{�i�<yV�T.d���a�h��x��o�r�'�@��ET�:k �C��ݎ?��	��Sb�m30F^�I��x�A�\z�-#ƛ7 d��ʤ+M����g�3��O`�E��b�`�H13�`��>O�H�f�4T1�<S�耴i�d��O�B�(2,�#Ҽ�˥��V�? �ѫ�̈́�^F,���hZxd�5��?	�H��ɷg
xh�2$B%VnA�T�]w��TC���O \J��5L0� '	ȵch@��C'Wd]�4c� q���˒�<P�A'�kL� +��D�~�oQ�-N4:��'T�h�ڔ�]�8�H��A�"�L"e�F�O�ȍ�sOT�`H�	NA%Q�d��L?�|^B�BEDW�Az��� N�c��G~"�*#�.��ǔu^9�O��4SG��J�ڀ%B�K����i3tת}��,@ ].��D�-�џ,��j^g�xlQ�N�	�(����)�d\	�"����)�	� ���@�#��y��cE�"#��c`o�<N&�3�	�&>TB�	wN�h�,��Iv�3EGC�R�ba���Z�!�
��6���	�S�f�]�z f��BL�%IX���7�Y�2C�ɧ<���b�	�j%�-!�e ��t��J/3� ��v�>E��'�&9�� Ю��DR��� b<�=K�'.��y�E��(|��M�Z^�-3�'Z���� Ô�ּ��ɉ��X1pd�.��u�𫉷�D���\G�Yh���Mk�"��W�6���,p|��`#D�<�ב^ɚ1b `��K�ި�s.<�tz��Ĥ�- ���|*�NT3Q��!���Q����dCs�<9#GS�!������rX�tk#,�2v8�I�!;H��ҧ���� p����F�*
�t���MC=�!�D߫ ��)5�H,�t�
U�,��D�P���� ���p=�SJՔ���:�AI�f%B����Mt8���#�5��n�c�~��2A4�uH�� ��C�	8?r|д&�& �I�pI��ud�"=)�E;<�}���T�K}�����,i��q2�I�'O�2oYi�O-����2�"�%�$@t���'����EC����`k��uP�mhsKI�[1�3H>a���OZ���σC�L"	��H�2�*T"O��`*�|ꭉ��ψ
��m�X/� �"%�ym���1��4�%eۧ��yræ�@]����	7MhȜ(����`�b��D��uX"m�:g6	�a�����dZ<{w�d
ד*'V,8���C_���`M߇Me4��>����f��`�4��C�0�@�BK�����~l�p����sBB�	I��C'ܥn}��"#ĳU9�����>s�U�Ot�KA	��wq⌳L�쀟w��� �i�1V!�l�,X�A�'$���*��z*��3��-��p����a���H��ē2N퓒τ�{��Ov���dA4"��*�0,u�����'�h�P&�O�Z����</��T����aH	�1+N�%���F[n�h���Zt���V�Kv01 ��'ᠩ�� �/k�Oj8��!�Y�$�I��H���2�6)p�ě����hd,�	uZh,ۀ�)M���5>h�у��w7 0�j$��� C��<�'�@��!�h:p�%>��;C&ht{Ɗ@�H����8[�`0�ȓ/��� E�}r)�r���aq:�l>�Hc5��/g_�Ӻ� ��p���&�Ǉ���R�_5Cw������y��۲f}�Y�qe��V{`��a�\k�)�ɥR�R��֩�Ƚ𩟑��CE�9�t���4��&�"�O��(v B8V�t4@奖�~�h����-#  )���V[`���� �O�ib4�ٴ0PwD�aw��h���:~�Yk�cG�/
�9q�X��)�8��-���'H@;�l���Py&D�n�8X�g�2D1r����+�M���@����b��F�S���@eN,���rFe��]2t�wh��,������8D��9B+�J�ǈ��P)����LU�&����)�t�l�X5"(J�L�g�'��b�銺h�.M��W'Z��l ӓh��dh��S,UV. "��	m�d1	�g.f�#!b-$��%��א&u��	�Zy��L�lT���-Q�~7�%����&|2聡!T�.��9���
9�a�/���U�q��L�r�ό�Ԓ�"O�a#�Q�T��abQ�(�D��'���5)�%�0�؂��~��>E�vj���yG�ݱ~\q0���e�4�h�,ظΐxR,�/.`I�Ql*.W,�8� W�^7N��W6�ֹ�҅��b]�+$taG{R�w+nTHz$c 
TH �u��ذ<���F�� �Ԡ����K�}�Q#��:0�D�#u�-�n���4#pa~Bh�;_f�*'L�&FU�)�U�K$��L��03v+הN��Q�C�Y�a���
���S s@�+�H�%ZD8�)��<X�C䉂. ���M�:;n�b@��*wư�2G�� �����(6R�"��:�3�$��mͦ9����H���E'�6�!�$[r�? J<��S(5�|1� �{Ja�b�!z*����p>�V�T�NX��PfG�<fE����i�KX�<a�N7z˄�C��V?qw HY �ċ��̸:��ԑ@�E�<�sm��V�@���;��� �AF�;���(��A�?֑?�b���i���{��؊M�`��3J/D�p`,U�5Lz���B�m ���'<���-����&>�X���a��&q��aC�ƶ}^��ȓg�����V��Թ��f�u��l#l�JaN	-/��@I�W)��%�ȓF�� �!���^�x9��ˈ,�~���1� (K���d��ظ@g3	���ȓ0r�8��9<�^�@��H�Q����#R爭h7�8�Ȗ^�t�ȓA�h[޻E�>�rA�մ&�\,�� 'x#sFZ%��Qb�-̳]J�=��L�8ܨ�m��q,�1
Ƣ�>�U��%�rt�HE�xY�I� +�.\�ȓm�6�ړ�`hpL��Xu���� $,s�]�A@��Ѵ{^2��ȓ/����kU'z�X=��Iֱ@h���w-n�bѡ�t��x�f� 
ۂĆȓh��*%���jV�	��A�J�}��~�=�Ek��.�$ �%�9PՐ�ȓ�B��"
P�y�U+����[�&=��.nD������X����;���Y]b�q���	6F����֘)�ȓX�.4�(0K���҄��
#*=�ȓq>��JQN��	���0ҏS�>)���3*8�"���%��m.m&���F%����F�
L���x3���NU�1�ȓ gΝBB��)���(r��D7�ȓ!W��B��#?T����H�L܇ȓ	<��y�]���
�B,Ն�>�0"
��4@�&@�l�ȓ.֐e���A.b�6	>J-���*\�Q�C�%/rhqq�L`��h�\���[�Ҁ�oB�
0��w���a�R;�ѳ��ȥdN@�ȓ��i��٩VeN"��ݮ*l$����LBVF̟yD
�� `<B ���ȓw�������>gb��� o���r�<�2���7ެ��'e��j�p$Gm�<�fJq�0�J�(��Y���\�<��S'j3��1!�ri�y�����I� I�ƣL̽Rߓv��Z0��
2&�����)��ff���ğ\"`ƭ��i�����|�%9��Q�����Z:����g�t���L��mzj�I��[�K�D-�ȓ~���c�M�7%򹘂 3�ؐ��8�DI�B��8�`E��±a8`��ȓ\)�� �ƛ=l�v��GhA,-"�̆��xL�*ϹX�����(RYf��ȓ:{cl�� ��Ŭf�p|��gA�(�U���Atj@�DS4}	�A��}r|�cG�X����ڱc��(w긄ȓ|Nt4 5���J	b�i����U�܇��l����O�T��b�m�Խ�ȓDL�m)��	�q{�E1�,��j���ȓJ%Q�'喉�F�P��\���q�ȓn\l�rI%>�(#
G�E[� �ȓ%mh�A�V+	���p�o�h�\�ȓNx�$�敲p������Ll3������E��	��H ,��CF��ȓea��Ek
�RNFq�0
P�u�Jԇ�S�? ʙj�F�o�hIcKp]#g"O�!� I�J "ԣvfJj�j}�"O�\�GP��Z�{���%=��� ""O*x{$2X�&�2�a�(���"O�@	�D�� �e��ْZS�%��"O^+tiJ�\^�j�n��:L �8"O��)u��-!�MY�M�"q�����"O�����ުl�̰���U��	Xs"O��PQ��.\�6��2���,e�"ON �	$[s�`K7o@-L"J���"Oz��.��X�vN�1o9��]�<�w$_���Yj����=��0V�<a�C:=���`(�
P.`h��G�<�2ꇣaИ�P�K��z"`SE�<�CΏhj��1�n������K�<�E�7b�x�*�Ǖ�4�j���G�<�%	@��:�#�,�p���E�<is�*M'��`�Z�{������<���3kN�PwD�;bT��B��z�<!��	t8��j�l̴(@�:5g�w�<y��0T����%.�����Kt�<	�hÒC��E��\1��p��L�r�<a&-�m�*���4(�j<ZWj�w�<1������5��#@���x�<�OU�Z�V��!D� )��ٰx�<!Q&�"y���k��
̙��o�H�<A���-0����Oӈr5��C�~�<I��S�u�x���z͠ �Sy�<�"�G4�`���އWp���Xv�<a�-ϭ<�UG<5P>]`pn�H�<!�吺qè�Ҵ*�9-��0��L�<�Я�!>)P����/ &|\�6��@�<aa��H:S`㙢i$J�J%lW�<�v�C9"G��A����`�"��桀y�<�c�:j4���yR|:���P~��#�0>�#)G7qD4���҅z�Ir��v�����jZܟ�V �L�d�éD�`pkg:D���ը>M� I�p���J#��
����)��}$2m����:^�`�o*!�̦b�����HW�c ���'�[�h�d^��d�"~J�	
�0��ι/���rhZ�y�%�_���AG-E�>�4�J�(���[�u0���	b��`x���1.h�X�gʠ �a~�eQ�HGR�Ǭ#t���a��/��a����yr�C�tFX��H�O����i#��O*$��ӭg<� ���M�z�0Hgɾv�B�	���Q�$m�1e��Q�@B�	�-@������r�|�򈚲2��B�	�"B�C��M�����ؑ`N�B�ɀT� i�q�^�hnH�qD�2~�B�I�Q��x@
G�_���� oN�l�B�<(p
��¯ֈU$�P��!t�C�#z_�89fm�(o���J()�B�I�|�dh�@.R$@�w�G
N�����FJ���I�o��0�o�"-�8 3ӣ^0|B䉝o�UB���i*�y����vH��=9���r��Q�[�ys2$�A!Sqp�)"�"OSeC`q��	��f| �u�ij�A� �T�\�c�_�"~n�}��}+��QO�0Z��{��B䉛|�D�� H�.	J)���Y>T�ΓoB�X���
��@�-�[�'�^���d�Uk��|0����X��!F�Ɠ7ި��(��v�)�����n���8 L�yh��'W\��ǩ�p�b=3�cE�s�`�;��N��ܤ����#�<0՟�$��dM  숉sH��뚨�y
� ���&��T�,���%���	�,����K���/`nPAAv�"~�I4S�eI�hSKX�U8S�ݵ<�C�1e��!P��b] `Q"j^;p��	)b��+�	&Ebf� Ab"O� ��M�N�֝pu����،"��'n����L	�1�^B"-�0!�D-�1h[I��ZE� @h��D,��q!��F�,+�m"dt^�b�*�	�~�@�T˝&ؚ(�v��Fܧ~�b
.3�&�)� �Q�$�ȓ2��9��^������ր@��*ń�\.hd�6��!
^��Q��~�J�D�n�BQÙ�}Ha�"��?�yc�2G<�{�(C�pR6d٢��<����'�2���-�&��<�߶]Z��$�ӄO�����a8�����G�6D����a4oXq��I�Nڼ=Z�fN�=hVC�	0LvL�cf�.c��"e�56ʞ"=Q�(F��}�O�(D	W+X�@���ru�'R����'\��9��©d�iH6��Hq����'ި�yF���YR�{��W�;E���N��C��$5]��:�-CVD��TnљB3C�I�l�r������9Q�,HŠ��-�C�5V���ʗ�M�59��s��N�BΰB�ɗ=�(�2�Y%��k�kL�E��B�	fD�)�3� (
�:�J-e��C�	bL�݈�(n%�#�f�ڐ�R��Oh<�C�X9-� p�dDV�yo�1S�Z�H����d��(Za��U�T�$�;1n�@0��ȓ5G}�u ��ֱ����m�,�'/ʍ#���S�d���Eb��P[�9�A��3"7(C�I�$<��!V�yEte��L�	��c�D���M[x�8�*�eT�1����a�h�@t8�,x*�0<l�	���K�
!0� *I����ƓA���@:40������u��ȓ\�dA����V*�����I�l�:���Mt��ZC��0q"	�F Jf��ȓe9�M�ad�f� ٴ��h���ɤY`S��ٰ�M�fMǦHw��:�ℒP��{B��p�<�È���"	I�/@>��dIe�'1��d�3;z#}��gSm� 'ɔ�(�҉�f&�[�<iPa�8r�nq)@�F$��5��G��֭c���������ە'�F���̼kSL�:V+�'�!��O�~��؉�k�$��4�jחF��č�L�v�2OLq؞H!�߀o�<�ɓ�10�z�r��7�O��iV˔�C�4�l��[��!��I4' ��u#˯u�B�P*�#��	���BqΈ~X�"<C
)�tr��Ә!X�L�Ș%q|rᓭ�W�B�6�<q��?'{:�H��#��H����'��3J<E��'q� �#��+ 6�S�/@M��
�'�������7Vn��#iZ2L��`ʙ'x(8��?����� �:��!1u�ԐTP0Ȁ�( '{"�|�w��O�ß J�N���R%h!i�61LY[��5D���U��(ul�Xp|�Ո%	(D�l��&K�94�E��M�6˨�!N&D�t"�핀�ȵɌ!rl��E�<��۾X�&%�0ˈ����Հ~�<��,�W�j��S�:�;W��^�<�����K`����%�|u�3-�\�<9'��
А��̚7"�Ę0&�CW�<����(�1��ݵm�^D�K�<9�Ė�y�*�k��BH��]1VB��4k,P��h�#+��ؙqŁ#F�R"?ぃC+>yr$*R����+�@�U�����?D��*7�I�]�E� �CK�V��C�>��.]�O�>�B"�����qd����t�2D���%�Ӑ0����R�Qwg�U1��0��&�ތ��I!d�n����S,�1pJ[>x����F���(�MK�6z�e �ꅸI"\<;�IƆ��x
� ���fBs9�pɀ�U��Vt�R��Ǧ���n�%4j�����3=M±S4�u�Fa���%�!�dwUlhIԏǘ�~�1��"A�6�8�Ň�@�h�	�^�(��Y�l�KN5wb� �l�I��4lO�mc���~�"��ZY���Z�Z�&���M���T)OhT��K�&1Kaz���	B@a2���L�<\�qoZ��'_|���I@��F�G2�'<\0r BvuJ c5�0J��,ZF�<��N���"L3r@p�:@�x2�K�	�q�Z�M#����a�� ��_.{̺]�Ï	;V}�b2D��I��̶`L�LA2��+�F�h��s�
����H���>F��/.l�		�� ��G��n��0��
��$^�u�X|�@bբ<3��`!Ɛ?B�!��<'u���u�C�N&��2'�9�!�$��y�0�+VS��x���-�
F�!�d�Z��+�̍u�6p��V�!��\�v��ѸCÝ	��Y k+w�!�6�.�����n��)ɟ6�!��|�&���Ԡ|�`�AAC�G�!�$~LlPS�%C�J�s���)L�!�d3 bлP�٫=����EJ�!!���Q:�A�䋯t	z��)S$g!�$V�/�ft
�mS�Z�3��͡XX!�D�t֖�:%L<�*�#�JY~�!��(>�H�'�Wf�\�j�)�!�Djq��[i�4�k���4�!��ьk$�8YE䒷�8�z�n&�!�DD#�,yaAʱ��@�CQU:!�I�m�ޅ��ș�jw
��@�ת0!�$�%OX䉡0�>e�v8�F*��	!�yh`�u��y������̘wgPB�	��Ș�I�N0�q"�)`�:B�I�d&,�#o<�����@��PC䉟�AC��%Kʐ�1ӅӏW�*C�I�.�:x@����Zm��K^�r�C�-m�bP��� (Dta[�n]�ZuC��,p�Dzv �%��Ӣ�/��B������ۃ'�����*o��C�	 U�mb�ʟ=.�2��(�#�$C�	�b���Xl�V.A9�,�C䉔����(W��A���R���B�	6Fk�����v��m(�A�H��B�%G�Y�a�
$�X�yp�I�B�I
[��Cl�A�m��iٖ_��C�IZ$�	c悱2 ���`x�)Z�'ɪpoP T�� q����_�X��'��%�dn؏"{����ķH5�M��'7�ZOܘk��%�dEN/��!�'���Rh˟x
Z5yׯݷ!���'��D8��J6�^t�aA0b ��'�:��"��A��8k!A�o�x9�'���q�I9����h��y��T��'ѢYSA�Kܵpg�Ms�p��
�'uX�YrJ� zG�	�'�ܣ8�Q+�'�� R��e|T2�6H��P�'��u���H��1i�c�'��I��'�4�T&�7��Y�o�D��'�d-�a�L/^�X�R3N��t-	�'��Y*R+R>>Y�A3>�$Y��'�ƤK�Qr 5�G��5F�5�
�'>]�#��/�.�����,]�6��'�FQ ��#���䘪S��H��'��E���?����M@Gې��	�'� q�iC�H٘���ዸ>�.�)	�'1ZD���K�CW��*� Ǖ)p������ VD�� e������><�a�"O��G#�)p��ha�$N9&�x�"Obt��N�9E���0D"^`""O�@����Q"t C�w�(�"O�lR���K�Q��OS=P��2*O��`aW�(�×�s}Bu��'If�k�nˤ/T8U��Ț�o`0E��'{�h�wS	E�E��@͕3Y��	�'�P�����
x������'�H�a	�'���z��Cc�>��T`߮�Ν��'�m�׎Y���4I{���'�($��]t���y����>jJ���'�<)c���*zh�p���ny�$y�'���sI�Z�2�.e�,��	�'2F Y����!{ć(a�4��	�'x��CÊ0U�L��n��%��'h��/YO��0��U�l$�'��p�c�R&��(�n��&���'1� `(I5j<���C�nb��'�q������bN�\�{�'-�DzQ�X�A��}���+\�n���'��!�"ƈ*�D���OS3 �����'�ЛA� �9��ɳ�H�aD��@�'^d��+���L	V�"���'Ji�m� <��p�B�<I7iS�'@�(ۢQq�q�Q$��F��X��'�!�˃0mk4U�WhT-<����'�"�H2 M�Ln�Hw/>:/R��'����
�m	�ٶč�ϒeh�'�p���*&�&���`A����	�'r�|T���>�l(z ΍7�u�
�'���pL��R�:4q�T��C
�'t�P�W΃�B9(�a�jT*�H}��'�y9 ��O�ި.�! R�M��y�B#�Mʶ�ɠJz`��U��y�ӵ���`$g߷|ˀ�b郟�yB�����C�˪v���
�<�yR��2xU�
3�V�9�^m��˟��y�(M�V�^k�Û�fL���'�yB�M9]U�|!���4�`]PWJ�y"�W3�p�u��.�I o҇�yBI��m�@����#�إۀ�ʨ�y,�(�
M���Y��V��aP�y���t��*��̕�^�X6��&�y�����As�$���i�U�%�yr��cj�QED�(}�`��ƥ�yү I� �;!��n�4@��y"�E>�$H�Rnѿr���a���y"m�$ހ���L�n����p�M�yr�ߕ%�v��" �2]�5{��@$�y�@b{ ���&v�����yҍ� �����N�R�O�H-���]F��rMآg��%���-�ޝ��K���z3�#<���+��u��}�ȓx�m�t䙥^;���b��l����~IP�
V/ɢ)���Q�Y���ȓx ��:E���1����'�|��%��`��8G�Ǝ|�	�a�4e�	��$A��F�ܫ)dx��Ȇ6.��ȅ��XH�r�C/Zb���!�T�C�|<�ȓkv��KȦN�e��&��ȓ2r��Kp�M`�v|�&ᑈ:,t��}�t���5+t@��&�zB4q��=�`�P�"q"�R���|_lB�)� x8�ԃ�<M�.=�b���50a�''�DK�}��	6oЍPa�� �u!�Q�>j�Ȩ2\�|��5!���喁B����VT�jVX��!�d_�f��U�_T�����Ԯ�!��P����5j���!K��~�!�&I"`<� @�4R� 4/�!i!��Ֆ��փЁ_G��آ��#F!�D�#Xh�����5�(@"S�țH�!��{��P��C��D6�P��"O�E��3|Rrd� ~44X�"O8���5d��	y�Q�Yx�Y"O�ə�H��	�s �.��,�V"O���s$�
#0fCwES���a �"OV��u�G7Y�b����P�7���7"O����%�&x@rL+��V�,��X�"O�P��ÂM��8����,�`!�f"O��PG�X[r�A�A ��q�"O¡�G�@�|�Q�Q���t��p�B"O�P%g��~�`�*��$���3v"O�Ia�
�P��L��O�X�\i�A"O.���mCl,B �U8`axl�G"Ot��vA�'n����b��u&�D��"O>�DK�G���d�=jnUR�"O6���S9�$�['���>�4��"O�
�R(��!`�����E�!�$Mc�ܗ*m����׌̃l��`�'�P�3a�J�:%Zy3Fn�&o����'u�1��n&+ L���?7k�'TL�YoJ+
�Z���)���@�'K���A"h����(�h�0I[�'��!,�Jm�!�^����,D���BNY��Q��B��	�,|a�O D���`^*_�|#��F�V�Ju ��?D�82� ��\$Q*b�ɻy��q��M=D����b��,\t�#�`�����<D�4�H��3����&:��]�:D�d����&�n�*fcC�[Rl��-D��b�[�l����j�-��s%l-D�\`�y@�4����6|]<��2l,D��r�݆#��h��(~��(R�e>D�(H�O�~Δ�[3��J<�0HĦ:D�( F���E�9f|x�	-D��p��{����h	l\0Q*D����gD�r{R���OȔ_�����=D�` QJ�,��p���Ə_OؑA��;D��K��܍n`0ä���!�����7D�����~�Ju�֍n4n��ԫ"D�|zU�Y&�N)@�֦#�b�2� D�(�BG�Y �;�Ӷ}�t\��k D�(�5�xAz�AR42��:��+D�X���
�pV��� �e���0T�+D�(8�⋤1l�i����+ �����*O����oL*�}��9z'֌i�"O�!b�:@�L3&ّ[���("Or80�	����s�� ��(��"O�1��U�S�P�B���,�d=�D"O�HvY/{{p�3��)$iQa�"O��فL�
��y�� a"O�T����0��]S&׍Wӂ�j�"O0�p��F�1����ƞ�ĚI0"O��F�ق	��H��e��c���T"O�z��%& �16�_&[\���"O���M�� V	S��=�b"O� F���$��W;8z���9?�0�#r"O~��dL����ɧn݇j�t�Ҷ"O��[(��������Řq.	�"O`邒���fD������u��i"O�����v���C��rL��"O̱JB��i$�sgN%S�ą�W"O��G�"\kGX;(����"O�I����2v������=w��A"OR	�R�@��I�aȠN�\5	�"O��Q�
+�x쁢/�c{�e
"OzT�!�	p�^����\�?P`tI�"O��apdHu�#хL�Q��"O�9�K�0Vc:�s���\�t�"O�����r~<���7Vp�a
d"O�P�@���d0�E�f\a��"O*Ia���-&�� b�!���w"O��7�ߋF�!8��\).�̈0�"On�S��Rq>`ڦn�:�1K6"O��rj�d�X��lʟ18�Z$"O6P
�-�J���!��ɤ%4�	��"OZ j '�l���	�u����q"O�|4��v�J�瓔C�"Y"�"O0 S�͘ ��b6���s"O8G��]����s�M�&�8"O:�h�L�6:��aš ����"O�xK��-(��P&f��Xs�A×"O�L�w���L�`xc6NX�PUj`��"Of�ӵb�[�tA�T,�(	��0bB"O�嫥�_�������ŉ.!�!��		���8bcڷ�h�T��1"!�[0z1��ʳΐ6@ P�����B!�ٴn�BE�"j!�!`$�A�!�d]�Y&b�!�(�>	bE36���!�,4l|)��΂z��D�#cE�!�D�[�h	��-�f�ȉ����'�!�dBz���	7K�>p�phk+h�!�dώ����d�$aj�u��$A�<�!�$�z�����,�Y���N�Py"')%���h&b�)]md4c�P��y"��mVb�!E�K�I4
���啲�y���j��0*�lL?�L��Fˁ��yb���\v���%�%E B��K��y��]�]�n�r��Ik��;&&��y�žv�^=p&�JD�4����L��y�=gȵA�Kޤk*8I���&�yr�Ζq0U�`	]K�P�B���y��8����2�h�@���(3�y�ҍy��B��W
�Qr��K#�y�(I7`Y�Go�P����0�̶�y���NK$�"�a�25u(@K ,��y�JW=H�\	@��Ͼ,6���2(H�yrE8>�p訑%�2�i�qD	�y�� �o���K�OA�9�0�*+�yr��,��H�v�J�5N��g����yBѨ'�6Lk��Z���X�n�5�yB�AV�2ɂ�/]�Y���l��y2M� ``�h:�	���Ь��`V
�y�m�NJ��㫕�F�S�$��y2��?6�|b:.�aC�y�'Y2T��sC���H�*�E��y"��Z@��A��m��A���y���gy.��l�!;]H�	 �y�BT阝�B9Hք�DfĜ�yB�:I�I��Λ�G�ȕiW�D+�y
� ��S�JF�!)�Ѫa
�#�h��t"O&8C%ҭ'���{ei�O����a"O>��pA�%A� H����#@�v]`"O����]�B��I"�W�\����"O���n�=bF��!�%�#E��� t*O�2� ��K�0�*��9br=H�'i���D�V�Fw4<
r�O	i-���'����pDQʅ�˨0��+�y���*,��4�F з�f��GȚ�y�ťg�>�{���w}�x"��Q�y���@���u�ϏY8���@���ybD��n䰱�X�[�z����/�yi��g� e���(\�� ���ա�y�J0�L�� ��=<Nlh����y¦A��e%�-v��bɼ�yb��7 p�IV��(R>����yBm0
��تW�F��BQ���y��� �)�G�&����D7�y��S�7��:�*ǃ/m�sB���y"��fc�L���݆*��!"E��y��ܶ4���Q3C�,*����I��y�J�dP\-�#f]�s{p#F@ �y��
�u'��sgir�!�\��y��װ^�	eX17EJx̙�y�*�g@r�
�$C2X�
	㥋��yr-��3�X�+��[�G^|@5m��ybD� d4<�an�72�l��&Գ�y��D�� �$�R&�oc����'�n���M�6S�LPw�A����
�'�
!SR�B	?j1\	uF��'�����E�/O��Tf;�"(�ʓY��9�̀�,�*U2��P�=3"��ȓ�90��8RP�Yg �?h�N���DīG�Ղ55�|�gKX<����ȓ1(��ek7v�)�NS�_�8ل�(t��3צ"�x�I�i :m���1G�Taw�$_��5QU9ZT���x��$ڣ+t<E��I@�N��مȓ{�)["�:�He;So�'w��T��F�R=�� ��OvA�Cf�IA`M��j9�)J6�Z�\O�@E獬sk��ȓ)7����疹 �$(��A�0=<��{�:����ϩ �y���R�4q�ԇ�-[h�"�n�:#n�qc�ҟo�6�����=A�fĆT\��LO�v̈́ȓES�`c� p�> zt����D�ȓ	�@�3e⇑q������ռt38y��*C���q�Z�B@�3D�N�"	��x,-J�@��o�#�!�8���ȓeI,I�ƅ
;^��I"�ӟx�zH�ȓ2j̫��D�#<̤ao�nav��ʓ!/:q���*wY�h@�c؁GxjB䉭wr�k��"h{nl2&!�*
B䉅"�t�.֒0}�d�	 ��C�I�hK8��v�?;����$8kC��4��M�r�O$5�j]�1�Ȁp��B��-46d�3��.l��P��G�B�	�==���w�͓$� �X��W�C�IW���M+
��%Q�([��B䉜=�İZ�eBn�~�ڀ����B�Ƀ4Rr��4,�v|&�Y�� C��<X���j��'v��"B��|Q!�d�S��Tд��4pA2AA8!��O�ȴ-h�j��{�\�W��?8 !�� @�3�IO�[A�u�s�L� �0�U"O����� �vT�K��fŶ5J�"O��ɀ�6vl���i�@�<�I�"O�p��f2,f�f���w��!�"O��p5a0j?��(�?v���k@"O
�{�Ȁ�ܨ���B�J��`""Oڬ���H�%9�����PI���Ǟ>����A�g�^H*����7���@�c�/0��O~�=��|�a¯��������!'j�a4"OI�P-;4rp�K�d�6��""O�XZ�B�X y����c(=J7"Onp	��� 4Z�1�"�"O���ǁ�~�]�!f8=î�b�"O��J�,�`ؑ�e�*U�R5�V"O�qR��U��#��5��E�$"O�@����%,��m`���<����'"O 2���,���ܹ̺E8�"O
�bC@Q�J0�`m�0
�`�;�"O���1����,zQ�ú|�(7"O�Xc7ŗN`����,Ϭ+X�w"O�U*T"�>|�V|ᤋ��&D� �"O�5r��T%^���#��̣#��S5"O�89�c�(.b�(�d�X$3���J�"O()����56AZA	N�`"O���¡�?;&ERPO�~�h�c7"O�5A�[V�P���Uz���"O0�î�2)�dRP	p�ӗ"O��4�/-��SC�ݑcUzS"O�i��jĒe��%r��()�y�"O&��ä	4ݜe�1C\;I@D���"O���­�0T"Ɖ����w8,�bq"O�\�s㗑��"�F^�d��d��"O�)S���Daab+��ˊ��"OtuhC-�	������=��{"O"8'o�4z��Y��j��2d��"O��VBH�*� �����"O����� u�R��p�t����'"O~]�`�߶6 i�� ^0�1�"Oʐ����=@�u�H�)A��RE"Oȉ��.�*�*�۳u(��C��'Aw� ����$���t,= M�C�ɦʖ=��e� *`�`WM�.�C䉑�t�(�@Lly��bƻ8q���d�>YtȚk��T�2�C��\�2e��<�$�km�@�`�XEe��#��A�<q���V\���l˥e�F�S,�z�<I�	gN��2!��M����E��r�<aPh�Iz�2��Ł����nr�<т�M��y+�R�K~�1���Cj�<����>՞��RKؠ)�(D��*Vf�<YF�ΕL��p�c�^�F��Ad�<!k�.g��8�U��hS��R1H�f�<�ц��5+�U��֒p�b��W�e�<A�g_�B�<��͙=<N!I��d�<!r�Y� 5-C�!�: i�B��]�<I���\G�7�L91��dkEC�y�eV�{{�� ���$��5�s�6�y��Y�Y�vE���b|3kؚ�y��P:�̘7�P����R���>��O~��b��s���b�U�`x���"O���"��@D�����7YVp�BT"O��!�eK �
�Ӛ9,�"O&�s��%N�x���i�6���"Op5���g!�����/ `�`"O� Xq
�$��X�ThY��9R�:�aT"O!dƄD�|�&��"�"OP����	��t�[ �w����"O��`'�	��Bf%N�#���#"O-�v�8�`!H�AX;r¹�"O |��l��(�q�L�;H�4c�"O>}�GMY�~�*]��GֽZFnh�$"O�!�gG%hs��Yc�Ԉh;2��"O��7��~:r�(  �{2Z0BU"O2�g�tؚ����"|���"On��N\A\�Ȓ�`�	�E`"O4ٵ��\��@��Z����R�'��)&�HJc��\�.�ucFl@�($D��SW��dѢ}ô��o��+E� b��<�O{��ЀgOL]@�p�#�"W48$��'���@���)3͈�ە�G"V�Z�C�/�S��?�t͗�`�,-�`�ޒ]��Pj�C�<�"
R���g�*(���Lx�<��L�m�@"�S/j�r2E�Gq�<1խ05i��z��X?s�|�yᩔW�<!��Zqݺ��!�7nr��qAGR�<	�@�<o'6�p*DP��@��SR�<!�F�$��=k�!�a�x��M�<��ǄW�b]9�o[i`�����F�<�����`���TmL5��EL�<YP�
7U������}�N�U�WE�<Q��K!&Ёf�ܷx|�'EK�<! �S�W4dd2�L���Ͳ��En�<14 L3f��s����l��-i��Uj�<���Pe��0A�@)0��� �L�<!P@�/IVe+���1w�EF�<��],1Ƣ9ۗ�
�:�lZ�C�<��o�\�6��-�+"�x��!{�<��Τ(�h��j��&��9 �@x�<�G��O��"beKQ�0q�O�<�,Ŧ&�rQۇ_*i��	A@�C�<9�#R��Z�[�f���Q$�\'�y�l�=}"T@a#��-ݶ��6�Z�yb�
�u��L�d��h�Ʈ���yr'�0r�~03��OE~�8�霾�ybƀ4.�bQ !��U�hu� B���y�%PT�D�p�ۦ�qI+	�y2�Ml���w��!
Į-bpD8�y�j�m�@�X�P�@T�2F��y�k��m`����2��EZ�R��y2�	+g���@v��
��A4���yBkK�J1���������]*�y"H�5����X������y�O�����˴8͞0{���6�y��@-vb�UO�#2|���n��y�gA)yئ�SE�6j�:�������y� 
���(�hW�8�8��%I���yb��3k���n�
1`�4�L<�yR+ �sPL2|�r���y��	w��`� Ӻ�h8��T��y�,��^^(��R��ŨcK��y�j� �x	��"��<�m��� �y2��]�LY�`�G�n$��G����yBd˲����Ph/m�VT�7d׊�yƣW���ɓg��*8��I�y���:m�Dm�5�B m��aFF��y�ϓ\Hl�:(�/���2�C��yb��?�[s.�����ª�y���崡K�&�� p$���D[,�y
� �� 4*WTM Hƭ�0�$"OjU��,�N��`p�S�9g���"O�l�uo���
��Dc�?U��x"O�D��#�6zCP�;ޤ=2��"O��I���ίX&
�A�"O��(���J/:����2m
]q�"O앒`˛�<��Pxʌ���"O&]���P�	�P�q��k9v(��"O��z� .J��(U(G���e"O������8r͉i��'��pa"O
��u`�JL����[;aT���"O��hϞQ�\=Zd��
<La�"O�Y V�R�S��p���U��Z�"O����"�M(X����9����W"Of�����M�S�@ 0�5Q%"O��)ׁY������ڱy�<���"OnE!,߭
"XA!��ʒB�ؘ�yR�m��1�W�s��q��畜�y��]�H�ڱ呖]Y�\����y$�Wmf� r�>!/j]%bX��y��U��:W"!A´ӃhA��y«K�'�(��E� 1��83�B8�yb%C�*��5q�E��x�v�GP�y���<���[QZ<`z���]��yr��MǸ,k��9n�����i�<�y"J�cB��i٢�:�O��y�DˊaΤ�!��N�9�K�0�yR�+3^�ԛ��^�(lx�º�y�I�*�<��f��\X�+�E��y"�U�hR�;��ÉTҼ���+��yr�Jg��S��KlRyȣ�0�y��Y i��(���W������y�C�%! ��qĐ CI$�f �!�y�!)�ޝ��� ����+L��yr C#k��QaAB	�v��p ����yJ� �8�o��f/�aV#Ր�yƞ+����T(��1���O��yB��
.���݉!�d����ߒ�y�愋vȾ��fL	�Ⱥt&��y���2�D%�7�rt+N'�y�I?.H`�'�­���A��y�ϋ��	���o��۵ K��y�Ƌ���zP�E	���ar��"�y�4-YLq���N>��`\2�y�˟g�Z`ɗ�F�F�J��"�yrL�n4��"�B,o��0a4l��y��nv��C�eM� l��C�
��y�I��[D �0Cӆ�t��@V��y"�͙��GI������(��yX0+BuaW�J8$�p��V ��y�U�(BR�q�f��&lܨ�y�	 �3_L��dL�&a�@Q�%ϓ/�y2m�3
�HQ��	U��X�6l?�y�ê�2�1х��If�	ض'N%�y��ѷ$4��j:*~�#��yRc]/4C� sdՕ˪q#R�X��ym�,08�Cu��2��*6���y'�8lT)3q�Q�ta�qv%���y�CH:�4)RqEΏ!�Xd��a�)�yr�
Q�m��B׷�с)U��yE�6���Y��K����O͌�y��)/�j������ l�yr=n��]
W	�YC�$K@�U��y�!PI��I���S`:�ŊX��y
� LШ��4�m��F���5(f"Ol�*�@N+GT@bǦ�,u��Ӕ"O����D�4��Is�C_,,s�sV"O 0���0":P�K���[��8�"Od�kB���[�GR<ST��J"O��B�(��"��܀Q�Q�X_.\ʡ"O��`��R�2�dā�+^S��s "O}�E-އ�, S%D�p�P"OJ�Sթ"I.r����M�;�� 9�"ON��&�O @�!kUD�$5���[C"Oʀ��B�b6���碘�`�Y"Of!�Fo� m�8y��M&f��@p!"O(D)�� (6� �ύ"k�L(�"O(9�%���eX���nV�4j  �2"O�H(gI�I0\�!cV�:��ey�"O�4)�;JÌ���Ώk��U�U"O��K�OՀWҤ�@�(����A"On����Md{1C�fP1�"O�k!eʔY`��!�!��l��"O@h+�MN�b�A�5"����"O����F��d�T�`�~�<E��"O�)W�P<{A�͚��̱s"O�����	��*�M�sĹ��4�(�x�eA"�J$�B)�-1���T��M) 嘪W	���,�h4�ȓ[i���%A���Խj��|"��ȓZ�r�
��G���ԩ��U� $JՆȓI�a%N[�����21@b=��#߈�jQ%�0 T.q��O�=�,Ʉ�D=��8�`P�-�.���e�8���OZ���D��-mˢ���
���3a�?,��k�L�9��	��VT�]�դW�5�������.���ȓ|Ɖ`�l͹o�)����̈́ȓ����a["m�6���PǺ���7Z�@�f�*ʪy��NA�Aڜ��ȓS���S&�0��柖>����h,�*�PH�])&��2'nu�ȓiJ+�Bԓy$u�'5��h�ȓ+� �4-W�'X��ui
�5��-�ȓZB"��K�;W�<PG��7�y�ȓJ��9��bLy{��'�'22��ȓXɌ�;&i�:8�<��$U=/U Ą�558(t��\�k�Q�Z���ȓtBr��V �&�T�+m�5g�9�ȓJ�"�9�f�4`@�k����Bżȇ�5e�౔�å6/�m�/ה#���Ҳ�A�#Z&V��z�O5y"̇�]� �IW �|Y��*b:e뎀��a��,�K�D:�O��`�ȓR���恌.o�f����M �~A��oUb	 �G-<�!��o�6؈�ȓKV��vOȣ�XP�%F�\�$$��.�ށ��Q3����&¢yk 1�ȓy�LhB��+�Y�ӊߠ*D>��8���a�ѣ(��i�;�~��ȓ)���0��)}a�(ك��u�T���k��\9$��)Ԥ���YU�ņ���;�	� ������"����ȓd�X�"4�o����5���Ȕ��
S̙��Ib���Rɘ�.���hآ�ɕA�"(�2*N�\@��ȓT]0�"eeY/ �T���+$%����\/��!�*:.S���BW�9��S�? \a2�H�!+`�եE;/�p�"O�pK�/K#.�µ�Aō�+��BA"O�� V˝&�,�$�eb-��"O}s��E�F�,N�>��;$"O<�KV〸X����d�{��"O$����x��'�W~r�"O��Y�F��0����aE�_2d"O|�':��y�dF�MNp���"O�� ��|r�HA���0d}�`"OD��P<yD�i�㏈-�"O҉�2�N-���U�V-G����"O��%@'!�:E�0�F�#/V�@f"O�aja\�aڸj�o,4��"O���Fe�jlz�;a��P��h�"O6,!��	�����'�1D8�Ä"O������&hej�"(�&�<x�3"O�ث�⅓<��s��I��]I�"O<��&�>U��
E�Ҳ3{J%a�"O��Y���
��9b�;�|�A"O~�(R�h��e0K�;o�$�"O������p�9�gׁw^�AZU"Oz�)�`�qipA�Y'c��!)�"O�uз	�:���y[؉3a�E�o�!�צ|��8��Spd���[�Q�!�͂Iڴ�C#A�6~|0����V�!�$@�x��bs�$J[`��fb
�5�!���n|�R�^�7^ʵh�L�!��Κ้ŋ	!�G��4�!�d�rZ`�oYԜ���Q�r�!�ح/��t�a�*I_6�@��<�!򤃛�$W��(��W�X�S�b��r�~$�W�D�GW�5�ƥ�	\e�ȓ~ڜa@��0[3&���W��݅ȓ1�vI	jۯ7�:�б������i� E��OD3lv4���[�zU�ȓVV��:c�ϫ"�J�R�Bي$�r��ȓk� |�pO��c��}z�U6��$�ȓ/H
U"Ga4�����ܭh0T���o$�A�@��0f(�2�ω#����hʶ-H�R?O��%Bg�Xc�؅�B����p�W,����K:]�vB��+:������$a4ř�O�#|�pB�	 F1`eLC0�����H�;ΨC�	7Z��<ٔ��%A�B�T�G�GP�B䉫�l�)��^[D��BB�M{�C�I�)d�&e*�,R�a
�i��C�	
$t�{"CD�"\�׀�;^/@B䉶'(�y�N�A�41'ҧ'�RB䉳�0 ��^XT,��AQ}�B�ɐ<��H��҇g��]�7��&RB䉻r�t�5�ܴa�>%��&<��C��c��yzU��  �9i����b�>C���<hQ���h.R��v���PB�	R���A�ʟE�Y��bB�ɀs��h
�͙e:�0��-�C�Ir��\����	f�����.�B��*�����c�2j8���F_�^B�	�1��#@�����F�%�TB�<;p~�s�o���cs�D8&B䉠0~8e�g'/#���F�f�C��$���I�ҷ�\XA�W4=��C�	:Z�D�pa��&ߘ�x6n�>��C�I'0oPM�G�FUO�!��/��X~B�	G�~d�7JTm)�(�� ,(�|B�)� &�qDo��$E�U�c�T�wE�Tj�"O (�� �@�p�b�
9V� "OE�Lv�~\�R�V.�U	�"O�@X H�?���
ƠVE��L�0"O`�K�b�-{��R��
�$��)��',�Od��B���o���M^�I�dpQ "O� K6��'#d��+��ɞ�6	�'"O̠yhG<-�(��M�`
<i3�"O�ݳ%D�3v�!àF�hPJ Ip"O�!:D��N����MΒs�tm��"Oމ��=�JX���0�`�U"OjLQ�T:q�`X��
��OC��"O����aTlF��6��2B
;�"O�TP��E�myfL��J���;"O����D�g�d����	����5D�h�ǈ%?n2��F��4!~���2D��r���L��`�C.]�!�5��A/D��ˆ�ǁF0ԝ8����.@�s�1D����}If!��Z�M�،)Q�/D�t�U�#����3GԤ����Eo/D��[���*4�Z	 �źfuV(i�%/D�L��S޾��@�C\���Sv/D�L��l�BY��&�S��'8D��iq�&#�f䅧o�.��'4D�TC��}��Y�+��vt�x׍=D��;�E�vY�MB��45i��sg��s��ryʟ4�����;�'�� v�3&��C�!�$V�qr��X\@��Z��1�!�Ɔz�z�{����!*��G�	�{L!�ԊU�H3�R�,~��!�!�ƕO["��L�^��{�O�6Q�!����)�KÔr��Vo�9g+!��n��EJ�NN!4�(���̂l
!�D�#?A�iA��?R��l�l�g!���g�A�um�9(��hՂe3!��	��T#�/c!����(!�ы.l���X5,B��Rh	�]t!�DQm.L����ׇRF:�1-ΪAb!��nLRc��'$�QA�T;QP!���K�lA�
Б4�`b NC�]�!�� �R$��-�jal�K7_a�!�$M��I���EB ���lʦ4�!��:G���w�J�'�Q���'!�$�p�<h�J�5Rm3��ǐ!�!򤘭P�{�#�6+<չԋH
�!�$�7`�2�(�	�R�[PJA�;�!��߬/�m���ΩOxv�W�V�fL�:�S�O�x�rf'XS�"tEʩ9� 8�
�'�rLbB��s0��p��U\]X��
�'�nQ"�h�t�	� P�v�	�'�Ĉ
Ո�u�^]*�B�4Xs���'�i�� ̈́))|���gB��qb�'�<��F.�JY�až=�s�'��Y����/9%���u�X?°is�'��8�A�G�4�hH��J��R�	�'t8��$.e|���bsȋ�"OR��B�(�HSd�;T��)�"O��h�3�(!�FJ4��"O^�X��jU�P�Y�R�V%A.!�ڛ������)VD-���.!�P�7�(�y虻,6��W��i%ax��'��O��A���y��a �J�ʌ2�'��O�����7s�������U!���"O�)��j�?)%����F�?�]�U"O� <�z&�ɮ02n��1%S�I�"OT�A c?�:<k��VQJx��"O�0b���\i�]P4?JYB	�4"O�X"3�M��iaRC̿��@V�-�Ş(��ݺ�Cү=��a�+H�F|����9r�� ��Y"�,��#��3�C䉮1�htu�V�C�$`R#oܯwG�B������U�)>���i��B�ɴ|�(�:R&�>p���d��8��B�ɦ
�L����юѢ灇U��B��j��%�a��찤)��3�"<����?�AФH�R�V��v��O����7�"LO⟼�Tmr���AӠȿCGpL���<D����!� n�8�b�@UJ؂�:D�����P�{���E�< I��%D�6�کO(���#�&���3b�^�<)�(�0jcg[�h'���q�<Y�o̳{�ZIwl�;S|�2D�R�<Q3��6Q|9��3��Ҷ��Q�<!����^D8p���f��+OI�<�d_<,�48'"Lg�� (a�Nk�<�����!��!펏C�R��5iGk�<	�E�h�m�m�ʒ3'��DC�� �2�$cׁ{�Th�UG�2�B��o��[+�o�,�R�a�i�hC�9p�]
��ܮN
���e��w,2C�		��;5FK�	·e�J7�B�/�y[ǉ�.Ajޜ��=P�|C�@X*DP��]�T"
m�q��tUvC�I"?�����aڅhr�LYd� ^C�	�d��1J�W[�)Ec�)y�LC�-u���r�M��Uܩ�č�9��#<9ϓ%fpɢ��#';���*ƹ,�$��,LPG�ʘBt�av	�_ND�ȓ~�b��I��N�0EI�JR�FZцȓpM◂�9�� u"N���\��1�V@�te���� wo���jņȓvEp� ч!�x��	,�ʽ�ȓIp^�� l̇7��p"W�g4^��ȓ'0��R!�{��A:6Fšc�Gx��)Z�(�,HoT���n��\�=�p�Om�<�S��C�^4���υܔ�*&ng�<i@��*��U�[ބ:Q	~�<!Nܢ:R���G�0u;NZS��R�<�d$̼s�0y�H,*��pá�Q�<1A!��@tvm��L�G����,�N�<1��6�Tp������thr��R�<��Z�cPF0{U%�@��mPr�<��Ε/�Ⰲ��4�Z	�s�LW�<i�M�H^������a�eS�ɀj�<�OҤP�d��ƪh�jl9�#�o�<1�a��bܾ4��)��%6.HQ�
�o��$�'�H�@u�� �Ht�J\2p��+�'Z��h�
0�Z<hBe��h�1�'��p��LM=������?rs~���'�t)����8�Q)��ӱ_�@`��'[�8�aʲ0!��K��l=}3q�<D��¤�k���@�Bw��}�0�-D��s�gS�{ì����N�ڀ馅1��hO���l�� A��[ p������n{�C�IH%\<�`�I Z@5��5N@B䉁f����)�5H��T��\�4B�I�o�$M	�鄩jv��AT�[�N1�C�	.:� UX�̡MX�(�EY
��C�)�  XZ�b�j��`
��1|���"O���oM�(�)#g� D(S��Q�O�,��ukD'��)�e�zG����'��w��Q}|��%H�u:����'��0`X,J�6ii�o48=:�p�'��x)�PGw"��#@�5�J\�':R��Ԣ�Q_��#sE��,�f��	�'��B��E�)RII���	�<m+
�'6R�j�Ւwb\|/L�x��I���'ўb>�v��R����B�^�bD(�r��t���I� ��C�_/�ƍ�j�3�RC�Ɏ+��	S��C;V�q��M�Yk���d^���'�84��s�0��J���<��'��v6Yo�AB,8Aӎ؂�'��KއFXn ���UlP�����y2j���$Pq�E��(�!���_���M�)§��Ӏ>��-(7���/�
U�׫ ���HE{ʟ��*#萰_-|�+�L�75R����"O ��4�#�6�Q�N@���')�O��@��i;4d�P�O�B$�A�"O0�S�h�=)$Tݢ&
E�d�е�V"Oj���(ьx�t5٤HA8ʪ鱶"O.Q���[��}����"y�a"OL��	X)FԠ��fƷL�F�A"O8�Ra������|�~4z1"Ot"fB�	X���V��=ps�7�Ş	U�� ݏ&��+�9zx�ȓi�$�S4(
�h�r���%�XA�ȓD���[��Y_c#
6�E�ȓV  ��J�!��
"��e�	�ȓ:}B�ʓ΋+TC�8
���=�p�ȓ��{f�ԁol��I���u�x�ȓ72�
� O�$����Ń�GfՅȓ8 �P7 �>�� ¨<(�4�ȓ9b0�����0���ĊL�o��Ňȓz�tze�;P�X< W�� 7�FP�ȓ ���`�AH���a��I��l�ȓY�p
�e�.tW�y�A	N�0,�Gx��'9d����ZB��e�^� �Ρ��'�NL��%�*w�8;���%O��[�'�X�&U�"��X�3� E-<�C�'>��������M:g�a�'���� $�H�vn�/,��'�0��i��N���+�`G�.� �I�'8����/���Ҽ��cH�"82q�
�'�ʘ�W#�Lt��uDU!����	�'��Iբ��[_�يŬՐ�,4��'�����.W+N����� jyt$X�'/���Á2OEԽ�*�f�F��'ƒ8R�!�m�YY1��[����'0�!c�:�j]ȁ/��LPЉ�	�'��d�$AI�}&,(qa�@�=b���'x6mhfW4 ��Z�' �<��5�'
���T1R���oH�!!6=(�'� $�V���?g�Ē���fF*L�'�݋P�����$��d���'��HdC�&�T�K�$�R���',��y�K)U��!���X M�T��'n��V�S�kC��RjF2X���O��d?|Ore�SB�+��D󪀹\'x��e"O:�ٓKSp��YtHCW/4��w"O*����YJ����@�q��"O�UzU�>s����GgP�1��"O,����('i�X��ŋ�'y����"O� ��L�Gb��
� qH�ѻ�"O:������/C.�� Ȟ -\<;�"O���P,P7GL�����+h��P"O�`�e`�z�B�[e�W)0ғ�|F{���Zh6��QV��`Wz쫳cU�6�!�M6 ���������8Rc�y�!���i��tsc��8�T���D�	{�!�d�!*�DɂE��5���:!#����'ўb>��PKи3nq�� HK4[A�3���<�'�,h��26"� J X�S-NZ�<1U�/,,��s�3!�ѓ`�T�<��A�W݆QK� �z�nQK��O�<�(L�g���,�w]b�
��I�<����W��[5ÍvG��Q�^�<�P�Y�n[�@�E.��sv��<����ӵ���{g���>s4�r�
=A�B�ɝu��j���9iء��`��B�	�X�f,x�N&D�҅�Z�T��B�	�7ȑ��O�hӰ�j���'	DpB�	=$,\ !�N���wA�~��C�	:*� F��_5��@���3��B�	�/�8"��ӥHtU��j��9��B��ퟠ��A��ଃVo��J��A�#D���խ�z��U��W0\  M��"&D�4�&g�/-�a�� �+X���:D��2�%4�8їm�.�
���-D��Ԅ��h�l ���J���H��y"iD5���� ��8#�$~��
�'��9Ђ�\1
~�I#��3=P ��
�'�Dh�RЋ��L# �+b`�O�%	�`�7�
���N �1�"O A���� ��� ��B���"O�a��	��)�֩���֧*ǆ�+F"O&�P���ھ�;��,I�>���"Ov�br�G-@��(C��jB�"O�%���� .����ϋ��4@"O�ᢅ�0u�<�1p.ƒ|���3"O���i�4����K Z�*�"O�1�䨊T���ѐ(�9���JV"O,�S��?N,��$�3��e"OnH���L�u�8cǓo�Di��"O����=찊�#C�&��)�"O~�p4��1#�aMַ�X�0�"O��[��%;�3�E�4���pQ"O>]Y���R�$���0A�h���"O�A��/K�Bd���D_&Z�����"Ol�1́	c���P�F3Bx��"ObU!��߀s�rɲ�#�	o�p)�"O�}�'�)�!p���9e�]!�"ON	�	ՈwhPa4@A�G
�  �7��|���ȯ"��H9͂�dtѲ�C,6B�8��	�DUP��@#�����Y/A�B��#B2�0�ѪSQ��}�#�lB�ɑW�"���y��1)���2�RB�	�A7T<r��:�����ę�
� B�ɫZ���e��h�>`C�-�0T8PC�	�K�r���( ��Iؕi�BC���,*pL�)�D��ӎx?
y��2D�\������+� i�L��-D� @u��U�(�Æ(O�9Y�D���+D�0��/��^��݀�(ʱ@}�$*R�(�O��c"��`k�,p�Y�h�cѼ��ȓy���[�#VA�ą6�p@��E�|����	5����D]?=X��D|��'$�>� H�yv'H�F"b����{�<`�"OH����o�4I���u��iR&"ONY#s�L>m:~d�@�� �~��q"O���#��>����)X�����O��$ɸ;����
�c���r�!򄃏k&�!��Ðk�:���#�9%�!�䚏n<p;S-Z7�P��L�����6s>Y�D
gG(�E����yBH�K��#�隲aZ��I�m��y"��5�=s�Kӭa���h
1�y��2\9��{T�Y�^�����y�%���,�C8"�� &�
�y��G7iü�����'��Q���
�y��=�*d��;i�4kGƸ�y2K2%�� �̆7Y}���mޙ�y��tW����'<�L�����y�b�z����D�:��#�Ƀ���'>ўb>! G�Bz���1(��Z�ցp��=D�0!��6kne�NZ8F�`�)!�7D� ���VVpƮV��8��5D�����ǫy�4�S�T',fXhB.�O�ʓ��	
&ğ�#��ٗA\�em,���!Iz!�3�!l������YL���#���!��@���
�ҨK�>��ȓ���'��� |1J��rx ��~n�1I�H�V�<MIq� �fX ��%eI�0R��D�7
� ����<uɺ��8}��h��A6fL��	Ay"�'<����ߩ}����(0Kq�	�'��������"s@�q$Y$��y�'�ȅ��b�~�:�7o ����'#���L�"�Ղ���~9~k�'~D|��@Lzcډ����w����'|1����0|4��rF�v�j�'{R@چ#�Jt��yv�M�C�h�H��?���?AƁ�7p�0�H���"8����UC�'rў�'Z0�Ĥ�|���娄d�Ja�ȓ1����B�Z�k��
-� Ex��i>��	�S�"x i�!QtPջ�ðj��B�Iw6V��q͑�9z:q!dݏϞC�	j����g��R�����Y��C�I�4���P2���wZΈ�E&:`H�C�v5T@�l�d�h��jC䉮:i�7ߵ �P����8opz����4��P�mX6�j�dI���)�.*�O��/���3U�2D��m�%:��܄�*���H�ˆ2Xz���CdM$O�x�ȓ_@�Җ�� ଜ �bG7���������΀1+����F�t��4��e�Z�p�@ ��dc���/ly�؇�C�wS�d#`�q��Հ��
�o���qbH�[�F9]��$mĺN��T�<	���i��A�B��S�9XE��I��LZ�!�D
/D(䅲��?BT��U�51!���Y��}I�D(=̱1рl�!��G�18P2#Ι�V9|esR��jU!�P�f\� Bw���0|���EB�p�!�!��m�ቁ~fЬ��o�!�_Jl�(��-|֜�$M1}�!���+\ɪ��p#ބ8_|�%�6!�ć)pJ�����hFr03���N�!�DB!+\�H����I?��:eo�9s�!��J<uܝ����:"h1@��_ ,~!�DI-d@N}:����*H�u��O�� Hp��.�/5x�	��1w����"O*�	�,Φ:t�KW�� o�U"O`����S,Zq�GJ];���"OƸ "��-�Hx��ȩ
�?�y"�$F*D�R	���7���y�I�!��us��=X��)R'���yr�R*!�>9X��-�
��q�"�0=����6}l���4�M�zT�j�@��y���+>� ��qO���c���$ �O���#Δu�}����JOf�h"O6����v��q����_F�)�"O�v��C�d"d
�Pa� ��"O�����C�؍�F`�0oX���"O8s� {Rn���
D��ȳ�"O"(��ŷ9�=d�ͨn��`#F( ��|�����'����Q�'b�t��GC_dTI
Ó�hO�i���o���(nK�6�x-@d"O���2�V�D�\��CGW8	VH�e"O�ق��RDfᘄ��5T�u{�"O��%�.t<aw�X[��88�"Ob%�3D�s�����3pZr� "O��2Q	�H�`����RK�}ʅ�'T�O��	DƎ�vX��D55��5"O�`ș�>�*b���/&}#��"|O"yy�d$f�qC/�;t�=��"O(-���'IZ,�t�#D��y��"O��*�E@�j�T����+n�>I;7��l�'��	
9�0�B�Чh��횄�\�0	�pD{�T�8�ʄ/�v���A֮�2��iu@��<9���ӶQ
<�IqO��W�f�����C�`"<a���?��7 �Gy|����������b�!D��`��<���!�O��ԡ#	!D���ЌD"'�Z���^1��=D� �@F؊G�H+�&2uR i>���	�mb�m��Ym�����O8i�����(�I+9�i�
YzР˷kL�0nC�	�p���d���:���g	�bP��	~��xxr(;������	�0�p�W x����	;{���#�kR:`�jL��Gů&�C�ɺeoV��g�!��*Ŗ7P��B��(W�@0KDbC:r���k��S���B������˃�*�5��<v��	{����N���F\c ���Ḳ��!a0"O>��de||4�P�&ɬ�r�"O��6`L�|T�j�b� zR?O���DB"
>��"JӠD��$�����
�'>��"1b�X��@q��ܧre }�	�',f���@K��9t���V��	�'�xz��65o��ul@�JJ��'�,-h'�o����t�	��)!�'<h��A��%Pb�,\*p%�L��y��)�S�08˕�R9$�K"l�?�2��e�I_y���YV$���0�>f܍�����!�T�6"&�#38��W*��!�DZ����x��P��	gK�!���l�4}�s��	./��2��`�!�[R����v��/Q#��[U�^(�f�=E��'Ɍ-�@95-�<��M�.5>�`
�'z���R�K� �Ѝ���F.�0�K��d3<OZ$r���_,X���k6ʥ"O��ѓj�1jJ���ᘍM�2r�"O��r̞�[tL���MؙSs����	x�'~:M �Ϝz� �4㏣%u>	�'��3ǁM�I��U���ߕ ���y�y��� �Tb&	�Nl�X�!A�3$�PК�ć��P�0Z���!=F�0�� v FC��"h��O-�XA�[y�NE+�'Bb���>+�@m�$	��_ ��'��x&��/���ιd � @�'�r�8#�Z�c.���I
��!�'�����12�Z��@���8M���)��<���<q�`�R4NօrE�0Çi�R��F{b�L7.�*��Ȗ�0݀�P��6�x�'D�$xQ�C+x��%- XJ���'����M�$%�T�WQ@H��'��d�Bb�X@�$fܹҒ�I�'��jF
�/w�ȃ3��3	}�3	���xU��J�C��h qf�P*l"Vчȓ+�tX�l��LIj��Z'e߆��'�}���??kt4�Tm�R@���4�yB��R�� V*�-b+�I��bG�y�!�*+Wl� o�Tu]A�$��y���<1gDTZ�G�H�F�ϵ�y�nR���5)��-S2d���^�0>9I>	0�'��@s `-"����<�I>�
�Mм
4jGF���mН>!v���h�r��Cl�1�����O�t`��ȓvk�ȵG%Lkr/	�~����.`8���"]�D�Z�h��U;1��]ʕ:e��&��##��p؈���V��$0򏝛\$���陨����	s��UU�Wꛌ_X61KǤT�O�x��y�IXLD�3�O_���`[2a�#q���d'��(_�R8�A�z;�xYg��w���|�IE����'>�A��,_0�j�seZ�!�䀣�'MD<�	Y+ z��F�|��Z�'�H���C�W�v��D	W�El��
�'a\U�GX��i��K%U �(z
�'66�J�%t�T�b�c�4#9�M��� �S���FiN5x����.ǚ���,�y�DiJ)`S�1+�z�[�%�3��'��{�kQ�;0ܡjP�M�BM D���yR�F	sԢp�gL�y�D��)S��y��S�t��5J%�p��q����1�0>iO>�r&Œ-���8sO�6�d��B��q�<�H�	?�]{uI�3yj
�Pҋ�n̓�hO�����)uf��֮B\�Ċ5��<	�*��+��-�d��:��P𒀘n�<��%҉2���e�z�.̓��o�<1��* �`�,����A��h�<�tI�mx��cCg�|*��d�<��Ӛk ��5M�|��u1Q��b�<aЩ��ؤ0b �0��y���d�<�Sd�{�Ġ���Zc��p�����x�jѓ�N�"f����(!��yB�6�d�qG�s�x=�ߔt�!���Z�aZ4�	�%��d�sυ�e�!�D[�u\�����Al ���4|�!�''�S�K��p��h�v�9!�$��PCr�\ ej����wa~�X���T�C�2u�s��,�"�;D��)���) ���\r� ��F/��蟾���e^�� �W� ��=(R"O�8{cT	fv���a��j�j�"OH�``�3f�89��K�/1�%��"O��ف�
���Nk&��"O��4��8����'
՝iall"""OR�1t����P�I%Y�f���"O� h8E�Y��p`�=��!�"O��xP&��}R�}�R�E3��dh�"O��3�OD�5��Rc��%S�F���"O�-�CcRh�p@I���C�|�@"OJ0e)��k����Ά��8p"O��XD��V]z���õ���a�"O|ȣU�ͭQV�(�L�.ϰ)*�"O\�G	?aL
7�OeHX*�"O�j"�.U�B�A�Z2����"O�	pѤ4QOY��蚀v�TU�S"O(-�@�T4�9#��W�3�v� �"O��%��8Խ�F���*�pȀ	�'��D���@W�ܫ���S3���' �\+�	'5�Ȅ�b�	���QJ�'	,�1�����X��=B02�'��Y�SH�?x9r��q��Ezhh�
�'i, KRhl�(\ ah�+f�l�3
�'D.a��g��7�^�S@�;d�.�a	�'E��
7�*Q���b
!+)�r�'�<t�P-�.
	;��_O���'���
J99�u��fR,І�rd̜§�#ɢY2B�ɱxS(���l��<��O�U�0�"�� vF4��E�Da�o�D.H�"�!u^���D�N �A�a�Д�4���_M�x��S��=qW�_5���k�G����Fj����*Ǯ!:�(����NU�Ѕ�zl��*����C�n% ��K�ͅ�=Ɯ����\��ѻ��t����"' �3�M�	D�,i��
mD�D��\����ʀ>2u�����np>���8�^�!�S2����HR= �ȓ*��Y�F�O$&�t��c�'\�=��N�P�;�V	3���t
S%Z�>��v�����L74O�)����9T�����	�ȁ��S�k^r�瘹v�����2�����Ͽ.Ѷ��1��6���ȓu�@�� �L����'�.����)&�x����${#�t���t䄇��b4R��c��̀�S�s>�ȓ؂ThFX�4"���D�h�����{�ܣ`�HL���M &���$�0��*�UCj-�.	;Lp��?�@x���Ch��b@�J�4L����0�le�3ǄN�^U��똀y@6a�ȓ P��䃝�4��Q�$й�^T�ȓP�^]��K�+>���Q��4cT`���9�8h�c��T��)��b�,g��؇ȓ_h�L�m�[ߚ����HEg����2p`t��%K�)����
��%��1��F=��37�4$��)���΁#10��	�=cc�K�b��B!�:M�i�ȓf8
U@@���k�<�4A3����}8ȵ�b��2�A��'M�BJ�`����"0&��eJ�#ѵdC���rV��!��oi�8ZR&�o��ՇȓE����D
$H�y�Ŏ1T ��T��L��ǟ5j���!� �-c��L���>q�Θ	���%�G�q<�=�ȓ?DAD�ћT�r��� �V���W.����]�d�!+W��J�dl�ȓwgl �p)��'���R�/]�Ml}��}pE��J���V ��<����ȓuB���7�WtjZq��R+JR���S�? �)feB"TDy@!�л��1ʅ"O�(�V��dl�d�ցYh/� a�"OZ��E�:���@@�K��('"O*x��ѡJ�E/��
�d���"O,E�e��4	��{�B�\0B�"Od$���Y�b4d�����V���U"OA�D�J&a2l��)��i�"O�5@啯/��(���O:���P�"O��0 ĉ$�^9SU'�M�|P7"O�	�%o�;�J�jBGB�A~�-p�"Oh��Ӄ�^�V�i 畼3����"O��x#
T���Cf]��F��"O�z?B���0�]k^��"O����d�t�\�T�I��txJ�"O�Xӕ��S�� �5�ߩh�h��"O�<���B2u	�`9 @�F�He�3"O,�ZaдJ��!��,�&ɲ"O�R����6���0��1�0���"O���t� �$#l)�CF6�Qt"O��C"�c܂���OT86�޹��"O �*��-EwP�y�(�1*�8@q�"O*� �o�!���!���R.p"�"O0ɐG���]����
��@ʡ"O��x�Č9�`�3�>v��`W"O|hQ2H��G���������5[%"O�h�&�#Y

Q�B��6��i�"O�����C�{ t}������jL�w"ONY�,Z<O��	���P�n4~��@"O���$%]r����fN�cN��u"O��@F�V�DT��o,3��[�"O�X�Ɂ�_�l��ՌO0�{T"O�h���ƬR��x��p�	>�y���S��ŀ%ʦW�xBwgI�yb�F9x:��`�RI���c"��yr(�ppi���#=� �"&��ybNY�LG,8�iǽ_i���f˒�y�HI#@O^�*��X�mI�]� �M��y"ċO����̅hUΝ����yRd�m�|�{�l�x�����ۋ�y"� |^�TP��N:WBl"�lX?�y��Ƙ_�(���9���J�I��y�NX�~$�Q[��E&*�(ɡ�c���y2`�  �l�a𠁡$5��26J[�yRD�2T���A��jY%CO��yb/��;�(��3V�Xg� DmG?�yR �,��	'�A^<p,�sc
�yR#$��I�d�ԛT���q�B��y¨�+$�8��DN�LҜds"���y"�� 8D�S&��
Bz�������yRW��a�@�R�L�:���y�+B�tQ��"��3G0@и֠�$�y�(A�f�m)�g��:/����A�!�y��ؗV�p�I��Ո/Vޠ:��V/�yblZ�L�aqFAT�HBg�^�<ye��>��0�f]�Z9^a��k�<A�`��/1 �`� ��'��;V�Q�<�r냘��	8�"�-cqJ�O�<w�)p�j(p��G�����O�<q� ����B�`
 ="��6��H�<9B�]|��`�cK� Ә(C@��K�<�TC�Y���Y�[�4�j��I�<ٰH�I�d� G������H�Y�<��GQ!j��p3���c�H0� R�<t�Q15M|�{d,#�6�Ham\O�<� �A���� ��*G�D9Yo$� �"O��@�	C�D���V�.0Te��"OVI$�J�=�$ �gF.#8��Q"O�U@`���$����%�Z>3E{�"O>����<wLE�'Ś(p�C "O�ٲI �%�� �#�ޫXmNYqR"Op�kI�c�>��v˘g�E�F"O8�'��?)�H���	d|I�"O�Py��޴�BC�4n��u�"O���''G��a�Ί-���!�"O����1R���%#��~��`U"O"�C%�҉@Ш	�A@�S���"O���%F�.�xq�g���z�c"O�m#w�	6J��t07 H/M�0dA"O��Yҁ	$� VL�Q|���p"O�����X�71��zV��c�Q�"O�E˂����U��;
c�ș#"OtX�SLײn��Ѷҩ
V$Y07"O.0*&(D$U���!�VN�qF"O�9�����8�OF�v���JE"O��p�� C�R�r�@ˣS�ĜS�"O❰���$Z^���s�x-��"O"XS�
) ��@���{[��'"O^��2A�:Q'��QEL]Oyp"OVdB�tA�4�!��*=�E�"O�y���=?�a��
�6��H�"O�9s��q���riA^'јv"O\�{����&5���!Q�5��8'"O�`
s�÷]0bw!YZ�9"O*=��蝲�(��Q�B�%�T�"�"O6y
��ʙ���#!��ڈq�"O���%P�-�z�rGk��Z�6`s"O��C1����U�7A�9K�05��"Oz��g�T ���h&��u�d0�E"O�<�SlI�*���)�߱���r�"O^E��:&��1��k�@��"O<T҆ŶQ|�(���Ů�3q"O��Mƞ%O�u���E��p��G"O�0��O�)���6�� Q�5�"O�E��mV�4�e��-H6��Q"O���t�^%V"�A���: G�<��"O*�#��L g��TP���,��Kw"O��0�'�kD<� !U�4)SE"O�Y�4��<-���B�o�H���s"O�qC�NQ�>���R�k@�Q�,iJ�"O�p�DƑ%��(8���?ofX��"O^q��Csm���D�U)P�,s�"Oܱ[U��	n���IG]0���b"O � ��A�МYR�^ \{$"O�$��T6tI���(����"O�Y ���wP��Pl�8D���""O�����A'$�ZdQFM�;Anfšs"O�������~�4�1Ё�.lf\��""O Y�ъ����-!�� |U��"O摲E��>)�� ��C���D"O ���"�0lL�9Z�f�q��B�"O��xB&V�=�����-d��{�"O��A"휛I
�"���6E� "OU��F�XИ��зv�B$�4"O��A��^cl0�[����B��x�"O���&�;%Ά����Z��m��"O���ȟ�7�z�!@;*��Q{�"O�M�pe�	(`D���	�/��EYd"O�17'~��r����I�F$s�"O� �	�O�_M�չG�ܫN�ܡ�"OV �g�(j���l�x�� �R"OT�a��,8�KA�R�`{�"O��ƀ�V�96�ՎdD���"O~y��a��kݠ��`�<v��� �"O& W��n�2�p�e�T�b�1�"Ovx�S=���0D�2ҲQb�"Oz����2=ެ�2���b`x�5"OЈ�獺P"$pu�P�M��"O
��䟓�4i@iG?f�K�"O�wOب=�T��'VVyp�"OQɷo)nx(��i��[R�y��"O��briJ')e(�&Jh[��+�"O���a�Ĥ|����P5$��&"Oq嬓��is���j��S"O>)c!�B�|���JO����B�"O���Ő)�(��7�Șxj`{ "O�]Y7-�)( ǈ�z[�`��"O~�sp"T�U�(`*U�W}V6�i�"ON�a�ق?�-��kN�:��@""O��`-ݞ+4xc� ݆%&b�C�"O�y��	�0P6E�ůBE�P�r"O��f�A5o��j7��U;&��q"O��	6��l�tUz�M�&,$�,��"O��q��OQHE��#�� "Or�@��,f�VIB�j�/d^ZEx"OH�٧.D0mmVM��^-\Ndܻ�"O6��U��r	�)HB�Fg����t"OV,��KY�Np6���f��
�"OF(�i?7~6�a�Ȑ07E D�'"Ox�!�T�*�"wN�\�2t�v"O�m�����r�tMQSσ1��)�v"O��	��D�[1.����U�<�.�r"O:��TGI5l4��"�
�6~8$��"O�̨VDS�q�]��Ƙ3z6�1�"Ol�0�k��=�d��Y{� Q�"Ox�yg�M�\��kRD�Eu��"�"O(Xzr�۟�Hi���̎tYZLx"OLh���ݏ:�|���!�{FT��"O��#_$��DPӂ�G\b���"O�ً�˃"~�2�k���+3cJ��V"O�T��+ �(D:�ŗrIx<("O��0���:=(���nQ�JLr��B"O��/����"��ía=�`�"OVX:4���f^Q�f�ƅ(�}@�"O� ���d��'W�"+^h��"Od��S�6��#�#�.E���H"OB�
�"�<(��(ǂJ7��I)`"O�ARu�E�B�QH0t��p*@"O�1 E�y�$XX��O�G��0�"OąA��W��a{�덬J?*=:�"O8��Ca�L�p媥
�'P��Y"OdPK�	ֿ?�� �
׍Bdz�"O�y�D��*�F�P�IڡZ�h���"O��	A8U�lp�Pg�;s��pju"O�#0���% E�y����"On��j̆�FuZS�T�ߒ�"O*��aP��V��1��U"O���U!r�`m���+}�
5�7"O^�Ԯ� N ��H|��S���y �&7+��8��ڐ9����'��yRF״��(#ԫ�24��Q�R��&�y�c���p�#���0p��e�R��y��E�kq�����U�"�� %E���y
� .yk �%0p0�t"J=��H��"OT9�S�=}��BQ�V[Q�`k�"O�H��L��]� ]8<̃V"O�0ٴ�W�mVf�Ή�}�F8��"Oy�!	�^$.q���/�F�0�"O<4��C�xE�I��4T��"O�����Ͱ4Q���ː2>���"OLE��ė��8H�)E/F����'"O$��<����G�@ؠ��"OT@Pbl�'{��Q��f�'��A"O4�F�|�v�k��
��%��"O��������VCQ��&��\Jd"OΡh�b�L<��޺p�4C"O��p��Ⱦw�1��� ��t�@"O��􏋨Y��X8q��"��Q�g"O���d�k��K�N%�ڡ�"O�X�V�X��y���F$C�j)3"O��KL�mw�l�បU#�q#R"O�a���D�gM�8�#D=pQ�"O�����ZB�|+&�N0_�ƨ� "OF��L�@���q�*ó?�ڵrD"O�1Btl��h��h��kӜ-R@"Oؘb�H	{��Uʱ�� +�m�A"Oh�@ <�D��o�a���"O��1��]�$�
A3�
�]�f�@B"O&,��)�*]�ځ���C�X���CW"O��CT'M�0�2��Dӕ*c��"O��x�G�_�j�9Q��{vr=��"O��9B��>
lP|2��+Z�P:#"O��
4^_��� r-R�q"OTQj���X�s���H�R`i�<�#"��`��	{�%"�����i�<�F�5t�H�e���,��Gc�o�<y7㕸i���b$�<���GPd�<i!�5q��lpE��b�X����k�<A�,ʂS�|�	B�B�&ƞd���j�<Q��O�h�Z����"���b�<q3D��*����<g�Ę��_�<%m�/R�p݃��@
9�v�PЈ�X�<�'⇠�j]�Rh�MA�Ux�SU�<Y����#$l<�)�N�<)�mʦ-PpS�M]N�]���d�<9���bΈ����D�D
<�"�_�<ie&�$�Ѡ5L�	k��$,]�<�B/ԘX+F=A*Ū	j]��$�X�<�a��iI�t��ҩ?�x!��k|�<�'ގ 8PHJ�k�$2R.�#S�M�<�&*�j�؇�_�E1����(Sd�<�`�"O�L]%���r��̐���d�<	���mV�I�7��wĀ��"	�`�<�B��<������9t�r���_�<9CDI.���:'n�Hȩ�#jI]�<!'o�=[�de�'�Q,��0�[�<I��B�nV$����h�V��K�m�<	� ��'�����Z��P	ԡBc�<A��"N�څڅ�9	��a�a�<Ip�������+- �M��R_�<���Ҍ1�`C�F�Rה�*�C�o�<!�" ���@*�Bɿ:����b�<q�%�������9d���+&�_�<�C��;R��t���ܵ;�@h�Du�<��iܟ:��t.E/x��|xLUX�<�U�P�f��x���M+y��T�]M�<ѳi�6=����]� �HIF�<� ����Ib5&X¥O&����"O�i:5�BI(�kH�r�0K"O��y���D�u��V9sё!"O`�H��)R[����Uw�5�`"O^�9f��&N��A��o4}�"O�%Ѡ�J!{+蔑���T�8�"OP�ks�V�)�e;Ge��EV,�v"O�����5siN������k�``�"O� �tIQ�DaPt�S�N�^���"Ox��的~��ePw���<�l("O�t:�.͜:��A۲A�oÎ	@�"O9��@�5:H���O���L�`"O.1�%��~>��O���N��6"O��u�ˋ:G�)�N��X�9�*Ot�A�'���)P)�-T��D;�'�"Q���h~���2�T�`$�t��'��Z��Սn7&e�3���D�����'�򱂇���c��Mj�T�/%8,��'t����A,u�1�2C�{0Tؠ
�'n�eCJ�����B��yL�h	
�'g�1IB0H��K�yqJ�	�'F�K�OF�Q����s���	�'2Hd���	][���-g$�9�'h"}�4�ݬE�T8�ph���!��'@���-�Z�2h���ϰ-��	�'dt�j�$�>sPR)0�Ω,����'`�,���<T^�����'A2���'p.�����L������<���A�'�m1��0{R�a
٭D���'�,�g \_<����&OM��pr	�'yV�󴊁g=���!�&JA��k	�'^�i1���)8rD�s�C!;�F���'��I ���?�>Z2��@�>�"�'-���0��a��)2��5���i�'6΍0d��-p������.��Mp
�'d�Dg�/:�t�`#]��z	�'><9a�B-p�~�y ˂�t��'�P�b�\YP�����i~^$y�'3:���\8Ŷc�'ج
%Ua�'�R����:% t���Lܨn�B��'G"ݒ��<@����7!�T�!
�'�T��R5f׊�`rAM�=�hl�	�'�l�8-ڭ&`8���-��&��
�'���JPN�� _�M��L�#9�1�'p.x��K���e����XJ
�'�P�viX�<�
���G� *�!	�'�z�V�J>HH�C��>T���''4`�4M������e� H��'�tY�1�>�5p��ΰ~�r�'+���i&�%���b,��'l����Ԓ�`+�B�X� �;
�'~���!�͓.���A7ȝ~��
�'i��;" �3'$N,ʁ��
yw~��	�'��$qR�W+_�j������nH�UJ	�'�<0�ηWڢ�js�C1s�P��'�:���k�s4La��7d��	�' 䜩�`�1/]�jE��s��+�'�*)e��Φ��Ĭ��rGdp��'�,���B�#&R�- �lڄm�$d�
�'�����G
N�K�R�h��P��i�<9�l@CD��o�a4@�Z��i�<�2��KT�Uv�;\؁�iHd�<�w������ɾp �U'�\�Ii���OyF=��딇.����?������ .�w�B �Z��FfQ�k[�j��	_��x�iV����L_�p�S ��y���>?�zMQ��߷% P�:��#2�X���'�a}2+'[����� �8�"��-�y��C����!�A	z� ��+L�y�cU�dT*!�X�1�
��TI��hO�'�"%��mh�H
A�3cU��0C�	K�"��Fk�����B��Q5n�,C�Ɋ\��2d��d�d(7aq�����n���J�$Bs��@�Ȕ�9^ �'�ld��	�/	BLse햓?�>ZƉ� �^��=}� (<�eK1��10W0qs5�е�yR�[a�|�fe�1sH�r$ݔ�y�ț�ڹ�v�K(m�x�X��E�yBJ��m&����`W�x�̈��y���L� ��E�"]ٰ�
�Bۆ��>O����	^L��4�Թa0=���+D�ԋ�
� �X�go�,����
*lO�����DW?8j�8�ͤ_ʥb�)'D�K5�Qsl�i�� wQ�rp'&�	J���'�^��U������OJ9��.�p���( ;�$) �M0u�h��ē�0=� �#������v�T=.԰���Cs �sG�������@\"!�X�ȓC�X1@X����E�S�|�Fx��)Z!aŎo:�	` Q�FJ���l�<I�OH�g��Lj�ɕ=M˾a�V%�M�<i��!E���I^e���3�E�<��@4:n�-�Ԏ�".��(���F�'Hў�'TZ�4��-3'6�j��hfC䉣8�R��E"υN;��30��@��hO�>2ɷ)Ӵ���mX��hQ �2��l�l�� �! E�/&`��˒�C7O���D��OIjty����XcdU=r!��@tL���󄒪`c�����]2W!�DU
 �1���؎CF��IW�בl��OȢ=�OP��[�o�:;�L�!���(	��:�"O���M	� wکq �(1CB�9�"O��AeYp>��V�6��p[r"O��u�5^�J� �+�9QdD,��"O���O�J�i�JL�M$�qC�-�S��y�-]'O��!�'b@'8RqR�Q?�yr�P�K�"���gR�^(���@/С�y2�.�Of�7cރu~�`Hr��F�6t��'��,�O|�
0ς
Z �U�F�\���ᕟ���)�O>��`"�O���q͘�.5���W�	`�'7��� �I���2X���A��oրB�ɜ{�xСE&�T��(��֌C�ɚv��Iqai��9Ӷ�p#�	6��B�I�f3����EU*��$1V/�L؆��ľ>���ҕJ	�l��ㅵ`��|�jLL�<E��6�HM�7%7e��b�F�<��iF�:��J�
Y2���f��wx��Dx"�ʚP�i.�
Ղ������*�S�O"d*�߀�&d�튞�t K>1����S�\=�s@�Ә*��bc��2��4}�΂`yJ|&���Ԭ�Ta�$ ��C��:$�̪�˪L�D�T &.Xv@���ѕo��$�,x��ᯙ)�L�b�|�Z�����#<��&��`Q�*�!��܃=�R�(�	�;*�� BV�	&�!�$�<`0�㊋S�~̈R@�k�!�D�"e���B�]�9�8�W�^�p�!�$ԙq���Ҁ�+����MT��Bx�� l�K6B�+U"��{׎hrD�'����<� hJ� �6o�Z)1� M d B�	�Y�$��s���5�*��I@�Qj�#=AQ.2}r��̞YJ6eB"G�!�h�26�9�!�d�tx��f�+� �Z�KL�0��)�'P��g��A@��c3e8�%�
�'ar	��G�q�c�5Y?|D�N��D{����ם+�B`ƄX�Qh�N���>��O�9���O�����-a�&0)�V�D��ڰ=����G�=����P�
E��jYx���I�<�2�ƹXO���1��9)�P� ��Q�<��lU�z�IDk�5�\=�O�H�<���5�ԑG��o����,�{�<�d����5�B,��"C*ࡓU~��(�S��G�0H���T?n�Ȑ1@��L�L��9���Y���/9)����ϝ�NlX!�=	ۓ��ٓV��w�*��kI�]Xj���x t�t�F3Ʀ��6i�����hO�>�ȇFEr<U( ��-O�L���J"������;��P3�@�@��Mˡ@������v�&�J���ȴ�ޖ&��i��h�,`��'a� �Crh�(�R��"O����G�zb���MU�^�
4�"O4h�Q�Y{��l,ƗY-�T�Q�$���F�D�B�9�"�a�04d�3we�-��D?��b8�;+:S�D�Ҋ��B��+b��O��d����OnU�,��'���f��7=�\`:�}4(@��TX�ܳ"�X2c�mp�K�'0*���'�:D�� ���6n,�@�'�"i�4�:S!8D�����֠:�9{6�^�\Y��1��Y��(O�b��bǡ��4����܇N���0�O��'q�)Cv*���P����Dwf�2��)�t`����2�%ׇ\����C�\���'K�M���"}:��	aK�x�!�@j�BD�gg�<�g�O	f�HU
F�T��*$��Y}2�'����,	)  �,ɶ��
&u���
�'H���b_�eeF�!(��K�١	�'�(�� ��/����-�.�d1��'=�dI�.ˆ.����k߆r��1�'������8t�4�
���WO�@��'8���g�ə*E�`9����M���:�'}@8qP*��J�RI��9S"�@�'&�
��G 5XPcs�&z�(�'���Faԥd�t�ӥNH�8���'�8�i�W $ɤ0�b3h��q��'Ųx����+|��rS�O���i�'~(��F�
I2 l�wjK�~�M��'���Kb�6'i��kB�Ӽw��d��'�6��@ګ*IB�����)w��}��'N��ه�ӭhɖ�CZ>|�l��'Sح�W!�&z.��0u����x��'����s�4-T�7��-P�-@�'�Ԅ���	;�X�@�/luP$��'�-r1'ڞl�X����f�n��',���D�
���4D߇J���'�Z�q�m��Kv��>�-H�'�BU9�'�oc�S�� +���A�'��ذ��O�x��е�'D|E�'k�	9�C�3��hҴ�P��fԘ�'s��qB��|�%����8Ċh��'���	1�8i�]A����e+�y8�'J`� 6L뺅ؓmD�]lhe�
�'��Y�&T�k�V0VB��&����	�'9�`9҅�r�'B�,�e�	��� 4u@��T�jSj�3���Qt�"�"O ���\*Q�XC[�ud���3"O��Xe����p�� >4���R"O������U�.`�F�2 FԹd"O�р&$ީ�JUb��X���"O�pK�8g<8�篅+lL�T"O����IC5D� 1�2-� k�"OFX(4���C���D��%g��C"O� ·O�"[)��)*�xl�Q"Of)J!��HА�1I�T+�"O�(���Ƚ\ľdc��=	f�h�"OZ躒�N�)/R�Jp��Н(�"Od���V
y�P۵���S�"O����=R��(wX&�Q�"O�50c FY��Q��T�^�Ҕ`�"O��˒���;� эQ���s��^?+��!��? ��d��"L�%ҷ�)b�庆�F0$(!�[�n�LI�-��j��M���� !�D�9�ݡ@eD��M��gд^!�D�;��ce��@h�I�� �!�$ݥ!IP�u���mW�����@�	K!�dЧ�Bh���ԬDQ�b�\!�$��8!�G�<i����E�>!�$W�*��l(��@�3i�CPo($U!�DS�&�BXi�F̯TB �5�+=N!�dO�:v8z���s�rd�����!��)I��rG�L�A!TS����!�$�?gDQI�hL�g0k7���!�D٭B�<��ә8&�Ȫ*�>5�!��1o8eY�DT+xG���*�
9J!�d��j>jeh j�<*(�&H��24!򤗉�U�ь��|?"ŋ�B��~'!���3L��#��O ��2��
=�!�d(-�P#���Z��y��@i�!�DO�q�j��T�j6���8�!���\J��Q�A 2�6ܺ�ڌU�!�DU������-��tp����ю;!�dʎ,G
�U&׷xd�VG�<<!�D�+�2���懆Fd��a��b*!�=yS ���A��1&���M58!�䊚F�|Y��Y�l�	���T!�[#��e�ૃ�#� ]�a"��8�!��84�q��G|�
��RI�!�ć1uY"�����&���×.M�!�DK�Vw>@� #��C�d�1EL�<�!�$K�YҊy11
�����RA�3X�!��8�[e].k~���ҫ�\p!�ʔ,��HȤ������7z!�dϳG�5�uc�7���'#�PZ!�$�����1׉]�$���aDۉp�!��		�0�p���h�<,ä%���!�$�/.:�x��dΆb��]��d
�E�!�$�o7����	j!NMZU Q!�DM:Fh�l2���&G�X1E ]=No!�D۠@�4X�SgDv�P�xw@\�FJ!��I�֦�Q5 V+v�!�/!�G�Pef<9ӳ9~`,*�+��<!��1�%��MIQ����&�!�DI	�
��@�Ή,Y�4XF�^;}!�ĎO�@�*WN�P z4��J�H!�F�B��ӅkYDF�[�	Oj!�$.U��B��ɩ^9�"g� !�dZ+7���R�(He�,�e��i!���6*���+��LS�(j
�HZ!�� T*S$�++ [��h�Tt1�"OD�ڄgM�^�:aZ�C�G�j�{�"Oz��q�Z3W�<�ib��8v�(��"O�9�3c�-_��]� 	P)n
"O=�a�E�`���j`� ��RQ�"O4�6O��^h���؍v� ��"O���E��l��
����t%��"O,`�X�_�T���&�'Ws���"O:a["�$BA�W�>s��{u"O��㌎�$���w���[���V"O��QKi�kq!Y;iQpՃ"O����Ʌ�x��&�ZK  �D"O�Y!傲` ����+���"O���B�,Xyz��"%lPD�"O�����S	p�ң����S"O�pXf�ۃ*��6m@w���J�%�O�}s@�֞�����������U�������.D�xAb U&�f�
�qz�y֬������BV>�k��'tѻ7��l����	�������$��N}rݫ7�D�b���b�b��})�iJ [�LB�2.�Dq� ���Sw7t�Tc���m��Wϲ�:�M�=%jh�}R�e�t� �*6�8. $����g�<�� F�c�4:"���x9�&��hƪ� �T�H���O�uF��O�a��çBŎ���ǣs���*��'�D�hT��~y��L����3����Eb�E�d��B�?ۨ ��-ޥT\"�I��"�`"ˉ�aS($�($]4��=Q4�ү�(�.O�\hp��)L�|�s@��+z��gF��:G�ԧF�xU3�"	�x�X�024O��_u���&H�>��}��eK���eg�l�.i�c��R�
T��_v���6��y�V@��|�0%N>N�<���-�'�p?��� 	YL%�VD������@�@�,�f]�mJ��
p�@�>�I"�̒<d�-�6D�����П��aPj!qL�ǵ6�TI<�C ��0)���0vf�"oMR�
��=q
�i%*�ZYz0!�+;���T垽	J�\�RO��J��bC��L]�ͻ�D.�!�J�8��.@�Y8�T��̓RL��R�o�� :�I��Ş�"�N�S�x�& �qn
-�T8���E !Y���D/N�ԕ�d�4B6:ҥ�K����@HF+v��	�%�FU:dȀh��px�BR]�%�EB���Ђ��G�.|���[�@Y.x��(m޵PU	>rJ�W�<�h1�Ot�;(D�L~���Ύ)�.�"fJ��Z�:DƇ�i����rM�/f�0�����Aap��KO�,�"�2�O|�I)	�q��
�/�����r�#>�p�A=h0�t�cD�9��(�`n�?�Ѥ�!Q=PQΰМ̊TCL)b	*��Q��$k�MȯM2�E�홇H��%� ��x2J�;"�ȥ�y��3��W�=$ޘ@��͹|�֤ލQ��lc��
�b<�1f��<�m�s)��!�"�"�cf����I�p	�G`J8%0�0����`3F%������CR��z�@y�U�`)ʇ�;!2�$��oe?^�W�"}
1iZ�9�n<�D�!D�"��$Q�JV}��H�Ѻ};����k����N�3{�|]y�M�7r{���v�
�d=��H��۪eח~�'W��	2�g
JT�6�Q�5�䠢��$ΐx��4{0B�7:���-��kS�T6� 	!s�ӱJ@~(;�O:6�Ji��Б0R4�t3q��?fÃZ7l��D��(N�\1�Do�ɔ)J�H�Do�(L�LѤD�c26���Y�m�,�8�b�U0Iaᆞ<u�1���(F:}j��� &raM؏�
��B�3�� 4V�hʄ]� N�(���ͻKF�j7i��X���	�̉�=�(Q�ȓSS12a�/r��a�$��$�P�(ue1%��ba�9}��9O��Ą՟4��{`ń�}Զ���"O�젤�V�i���b�*� )�=Oj���� X��דA��g��%�� �	W��@)��)N�6=x�
!d��(T �Lϸ�fσjR��� )D�D�0�� $ �S��6B`0R�&�G�L���IL�|j2`ފ}%���iY:+4$Z�D`�<�V��l����`S;%��YDc�4h1`���n�>	2ӧ����	`��t�Í�B�D���FԋX�!�dE6�X��ԾiN|�RQ�:���S-D�d���=�
R:b���wu�T��K?�O���i�./:7m�?H)�%0�˧,>�e��f��b�!�$�C�vɸ�`�@?�9�Ȭӑ�p��!a��>���#�kP<�
�g�-/���y� $9m����'�g�? Q�(�~�^�2s$�5n�r0��"Ol	R�gQ�b8�i�P��w�<!����w|�9��|��d8�# DO*� �'�3V�bM)n5D�T9�`�!EXq�4�� ep�DdA��(��I(ߓgS��[s�l�����L�Z�6���i�b��_�:�i��`Jl�c//X���{1&Йz�5�'�����"`��,���@L�\�V�x�+R�?�	��d�w��9M�O=����)v��V��&�;�G^&i��г"O@��ǟ�~�Z�GIW�ʼ���T:\~���gA>}�'[�r���Ç/B|�D���;bą�R�nHI0 hL��t��N�<�`V�]z���Κ�xh��"��Ɵ`#�e=��&���&�J,p�E�5�|"a�7G�`�c�gɊ$Lh��#з��=I�D	^�f$�6�O�� ��ޛL�4Qz��d<�S�lR��Ӱ&s����'�ZQ�GN�� ��� XY���}2@t�6-Z�^U�@-/�`MtjB<m%8��HC�'J�`p&�~����'�<#4���&�����W���P�O�@V�bJ<��n�f�� ��8�i}޹�W(_�x��)�1��;t�|ա�f'D�`�GHq�Cw��.��d�i���� ��g��m�K��s�Sg���4 ���"��67��)ӪZK��ȓ%I�Ui���ũ��ۧj3�5K��O2���O�i�u���s����H�O��A���jX����/7��}�F�5��$�4 :[��GC�cC��EL$����eP�Pya~B��KB��x�JH�d����hO�ѥbґt:ֽ"bb3�4��O6D)�ݖ!]4���Nw���'z�y���g�|x�I��D�\\���, ��a��
�4V���r	/�禅�C�FS�X[׃����h`e�4D��8pd� R�1d����k'�Ԉ@l U@�"E\�kA�ͼs�T�g�'Y��i��&�>�Q�ā^��	�A�� iH.U湨"��!T6ˀ�H� Tr������s��+�h٤��ex��j��[�a��� �/��Y.�����#� �[+��˱kïS���cj[
�ɕ"Jz����-50> ���,s=��R�N�y�i�00-yDU�jNrp@7-WF�xE0scБLL��$�p�nay����:k��,�;Z`dH��(��l��4��2'Y0���`�P�m��QC��pe#�T]����'V�B��pI�$R<��UEZ(|l� --�s��aD� o^xM�#��)�>L��I�B٨���ǉ�Vba�n�=5���(�E�T[��@�Y�AB
��#� \,�C��. 2��H	`���l!�:�%�$�gؿE<4EC�BC2		!l^"x��ɧ���N̢g[��k7��k~�4��"O���P��$9(��}U��x�c�<o�1[���B��)�E�!3���'|�X�پ��l2�K"/��'(�]��
<Uو�:b@�w$x"�)Z$��5�Y�!�|�^7V���`�H��C��+9�ay��#~�Hy��^�Vs���m^�I��ILoDB���7�!�M4qr��B$N����A�b]M��'���i���O��@G��)
��u�DH��`�^��y��Ù@z���EӫN7��נ[q�8���|�������3J^8%`�(sP|�'�vB�	�b�"\��玦L~l�D$ֆ h�C�	�p�(���\�0*�Ԫ�B�vB䉡�쨒w픈��QW"!.TB��:>�\h�7�_>o�d�	�%�*kxC�	�g�tV�u��@�Q�^�J���"ObQA��	�U[KL�T�D�P����yr���
� Ѐ�m>L��2�6�yBʄ_VR:��$ip�:�&�%�y���5]�8�`��7�H����y��C.Vu�X7!BY�]XT��(�yr�X'8
��Qe��\�8#c��y���F�N�b��*��Â��y2fP4.u�D�a��l�b4`i��y��Ǔ&s ��'�X�0Z�JԘ�y��>�,�{���X��[B�"�yb�ڊD�P�1�C��i6�U�p����y�{`%{!kP3eqę{U�:�y
� ���ٚ�he�R�^(�(��"O`�c��ԟ5�xaF�P�6����"O�(��h
#�T���N�=���"O|�:���Q8���FW��MP"O�`fW�=�*L/k8|)v��)�y�_55`�P���pgH�[f�L=�y��0Iq�ͳ$�=v�FC�ؚ�yR	�N���wk�;��[a�=�yB@L	!�� G�sFM��V#�y��+�=����o2��cn$�y�ɏ/�% �G��g�Rx9S%-�y!�M��J�>G{X8���y�o.n�YZT��;rPhj�MA��yB`�>��Y9�jNXh��k��0�yr	FO4����#"5� �V��y2a�	Q�B��!�y5.!2A��:�yR�,"|�h��vY0){T�ϵ�y#� ~T�A��.e��!�����Py� �%`�ڨR G��3��+�^m�<���(,���T�Q�J�V�ȀB�<���U�F!��aN��|X�[U�<9hT�W�d]zQ �f�>�
fM�Q�<9t@�n������ĹGٛ#��P�<Y����6�>�L\h(Fe�<���)\nP�q�\�4�@4�1l�j�<�R+p4�􎒣~Z4�c�[f�<����/R�@X�vE�99ʨs�![E�<��eYUt2��%�ސ@�l-Z�Ė@�<1�dݧNa�FXǰ�9�nGC�<��#��V�Τ؇䖵�L��B�x�<�7��[�V0`s慩?^hVOw�<1WO�M��@�K,tW���l�<I���c���
�H0,��C`�LR�<���V�x��ʐ:J�3a�L�<є�Z;�]��H�=�|�#���r�<QaC,)��O= ���R�$�:�'�f�
C N�}XK�n4��]�	�'�T��7���Kͼh�àԼ [�4!	�'����LM1M��!�C'L9
_`=��'��)Y�J�0:�� �be�+*0y��'fn�q�Ϳ;�x��FS�D٠�'/4���a�G_���r.�8���q�'8���$�V�w�ɂ�)�5(�|���'c���֤	O�`b@�Qq�81��'� ��g�Z��e�gm�&n�a �'B�ѱ%���I���~l܉��'.Xat������9�hh"�'��u���X\mX`yƅ��3e����'H�Rn[�Q���ȅ5)����'�*�FH�Lۆ����=dH��'h�0�ᜏ�����Z�Y�*���'uf�y���:�2Q0���oJd(�'�D��a�1=��,��mg�M��'�� �텳0��1���Ax1�'�~My'��ayzi�w��T{�T��';^�(%��=�A#�)N$\���'� PhE�Y:RJ�2��-O�ʕ2�'VV@(���U6����C�8��Z�'�5��k��)c�*>�0�q�'$���2e@6J�BH�����`�'�\�Bu蔔�t��vA�y�y
�'���Fdά]�@ׁ}�"���'�dY��?~R�Z`$S waA)�'�"�K � �v����;1ޱ)
��� �%����8��J)�B��"O�UH��C�Z^ D��d� ��(�$"Op�e�J{����Ab�6H�9�""O�9)��D:J��<�����M>���6"O{a�H�d�du)�ؓs.���"O�C��XVfh�%�߷` �(�U"O�m@Fa
�,4�<(�J�Դ:�"OF!S�� _����Ɠ%�03�"Ox� u�Fki�骄f]�8?<���"O��IvdD}��-#d%Ю7�A�"On���)U ]��2 0e"�"O\��g��2K��80�"�$2Mu"O�dk3��&@䭺�AU>A�ذA"O�Jv�W6@�z�pǃ��N�qr"Ofs�����\��@��
`�0Ӂ"Of�'D��l����/֋fP&ى""O:�Y!�)^tk$�D�n�˦"O�;4�5�ؙ���	�^l` �"O�d�4�ҴVܢP��ҚFs2X��"O*I�뚑�θ�be )Kzn��"O�Y!��Y5b�HhÆ�?��I�"O��Q LϰU'>��M
�d٣t"O��6��$0\�-��a��"O"���n��_�H��q�p�H(�"O�(A�X"e�%
Hb�U"O>D�B��N�`
�W5l���"O�@ch�]b���a�'T��W"O\�;�J�=B���"�1+vhÐ�'T�&�Ny��7fd���ȃ%E�g���y"�
C��YZ���(F���L�޸'
vI,*(r�@��IȄ�4�iҤ%�z1��}�!� �-0��1���j@!��`���b���?�&As�\9)����}�A� ��%24�@���.�p?�KZ�cE�A��-=X���M��}�RaئkB6l��q�T�J��|R�U.e���J�C�A,��A��@��O��ŬלX�Va�>"� ��Op�����e��0#T�Q��NP�yB�ѩ�JT��I�D[�O$N������^� �ɴW��l�DH����0�%N��}>E��O�TM���T�8 ��2&���-h��Z<9���I�^��dS�/[�ݳ C�% t��D��.{H8�rX�6>���[�,B�+��L��ҧ5�n�
JD`�I�R"�%;��4�0?a���r\Lx��޶U�|�� #�Z@3�2��E�ˆ�	>�:�`5��	ql��}�&����b΅M�~��UJL�'�n	�C�^�P�։�cIV��D�'}�~�b ^
k8��y��M�����O�XA��ΘH1x��I|�>��jY!C�bL*�FD�*�!�cL��<!��Ʀ7eP���	ѡ<̺	���6!5JS�#�+&�	ംV|�p��ɉ-6���B�'ؚ�ٷ��2D�����F�\�e�@���͏:B]`8I��\��u���b�]��.�W��Ʈ�Ge'	�L4pt�}�s��'�h����*�V��!ɸ��g��՛B�
d���;̚�x.ԠAH�,��))�	:V���6!���EN }ꑟ�X�P��H�1�,��.s��`����P�B|�⢂)M\�+����7���TQ��ƹY�џL+s/!%h$hx� s8$A	0�3���q=.U)�3��9��0�)Zy,�y���1
�ld�5Z @6|��P*��<n!�����%*��BG^���R 6ܸ�rCƚU��u36
Ԁ|���� 4�n(8�x 2��#J�agf�|(!��H=��� 3���F6�ͻD[�8�����
7��yL�"~Γ���e��k
y���3IH�ȓ��m��#��c@B��@ǌ�j4`ϓ>�qZƤũq���D�{�Ġ�r��9�0䳷��a|��_�� �UJ=S�< ���5`���v��4H��`�']H��U$�n^��x���
A�����dH0��K'�(��m� �w�(դ�;q������u�<�D!S�!hd@�T�i�l�G�ƱJ>EH"�`Jӧ����w���B��Ƅ�� �/�y"�	w&|M뒪ط[,��憣�yr���-��a��A��� ���d/S���a��Z%ApdyP6�'� ѹ��٩'#�fŝ]T�|8��ْg6 � �$�y��P�Njڴ�!� �|H��#=1�hߡ�֢}j�-֚Y6���mү`�p4�][�'�>�{��l�O�<dAK fuJ�:ԩ��G8���'�VYq �LS�!�(֍<�H5�2�Քz�L>���O�d���2�Q�=&P)�b"OR��2�W����I$vKh�i��iX��:��6P��5��C]�M���+�p!;p��60�����/���44��Q�IT�(�s4�G��z���� B���:���	1\O�1��(Z�**�ɗ@�X*q��d�IV��g ���'��A�ADrl#Bj{�Fl�j�f���	-�yB��i��:��gČ�I����X������!aJ�~�b�#Q��8CŒ�'�h睻c�. ��1E@b-��@Ƙ|��B��&�"�+dس`�p���j�x�B�B�cG�%�-7��qϚ<��[/��_>�K�+�t �@	�)�z<��	B8) ��ݎ,҈��}xV����@8������.?u�T��"I���<���F��EM�]�RTvNQ����#��n��'+ k�G�<�2���T�g��1�0Ɂ5b�zR��hh<���G�nEi2 �94mv��'�	?{"$PT�T�	#{�` 0h,*O�O%��ʴ�@���-�vN�ӧl��EI!�dȜ�B�XC��,�@!*��J"�����c���%�H���@�Hc�I����E�qAW�m�vY7�&O�(��vK"D��HTǗm�VL2�ǫ��	[WLC�E��+�% �ȐJ��ݰt�0�g�'ӈ�(LϠ1<\� �M�7kc<E��ka4Q�g�c�R�1�>faс�^��G���Q��k�3��MQ6g�:T��Kϩ+jqG{ҭL�hV��q���%���Sʪ|��/K�Ly�$ڮ1t9k�r�<Y��H�T�)��R s,N�zD�L�9�
�s�]: �D�P�X�)��s�P��!��&.Q��/�9�D�b"O$Y�ō���AN@Z���U�s�yЕb�8L�!��K�8x�r�g�'��,"��6^�Sw��h��Pӓ����H�j�~kE䐳+l����@��9��Ԡ��O�'EXl�b�J}��cႭq���kF�5�QMM`p%�0���Ojd��и�Ƥ\ ���,�d�b3��556T!2�u�8#c"O���!�6P(�(P2 _7~�d�T�IcE�#	��(cǑ�{B��>��CHO<�y��ٷ��h`�	|�`yX�߬��x�mC�\ؼ�C��UU�1����P|йu�J:A#����1}r�ıp%ǜXҨ�G{�dغnqbh��B %,���-Қ��<���H�F�RhzGE�%6.�c�M�0O���&�!	0H��u�(��d��qla~��n�X�1��(fS/���Q7,�PV��	 ��)ؒMZ�;���cB���ӚeX�q�'���
�i�%�*h�2"O�49���"F�i�F��-V����&"H�e���0B��l�X�r���k.���'"�i^�8A�e�q��8��Аx"'�0Ġ��@.YF�: J��M>�K�L˹dd��E�'�X!U�� ��!3� �w��m�˓%B21�3���e����'�h���AɟaOةؒ̍�8v����'Œ�kw�"y^����=0��msO>��S�2��ySw9�,�z#V�5*�(P��$� �ȓ-�$pr4-)y�&�)ъ�
4 ���
����4��E��O�lUO�� ~�5�s��07X� "O��h��M���1J�
H�"O���ծ=7dm0��$E�:\Y�"O\hC��Gt�A" �@���"O�%��x���`�B�!��A��"O�=J�	ИNM�0�$
� �NUh�"O���t��
���K��h�����"OP�)oL:h��@&�B���]��"O�%!��q��s���i�d�w"O�l� ���iwp �箚4C��;�"O��2����k1.���M�;���$"Oi�E�J&>�� b B��bL�Yt"Ov�����u�\!r�V^�İp"O���H� 8��`����/K.吠"O� t������(J�L1�D@�@Ob���"Od���ճbFe�1!#�YE"O�P�w+[�&�y�ؘ����t"O���KV�n�DA3͞	���I�"OHmp�D�Mf�͙�K�:a��m��"O��X��Mv�h�p�Glp|,�u"O�LR� � �>��È�sq�f"OV)"��&x�$���gը4t���S"O�)
!���!�ѡP{0�X�"On�BA�<p��.�?J}|�"On�FA�4h�0��^�d�B"O��y���/D5re�ȫ���!"OF����F�Z��U�'m�����"OiaTm��cr1��+��qks"O��@���|0,XK�ˆ
!���U"O���5_4Dl�I�W�\�܁(B"O����Nۣ14�0��uu|i�"OaZ���=0���%�o�t�"O��c�O�|k�=��N��D��q�"O"R�9�P᠗�^ XD�ʵ"OH�m�xӂ|�+V�
��@v"O60�C�I��P��v��k�"O�U�5B��*b^�@�/���� "Oi����ކ͛p&9�|��u�P%����?h��$��b���c���@aVx��� W!�ĀI9�dY�לp�>��?oB!����eK��Y��0PD�C!��Y�
Z�+��A�gr"E�_�g!�ċ��@`�£� a^�t�D#K�|V!�d�%��<�G,ľ9R�MA!,�+kE!��J����7CC�c�\�ڑ�K�s�!򤚧�X� �^���y�c���'��#<�����i:��<�c���W�Δp��:)���P']�<Y�lL5F��J>E��bW�90Ԏ�q�8� 4W)~e��A�1O�?�pb�7xL�2��׏� A��Œ%��b�P��E2�'����	�ҹK ���O�i��̕J��b�p 3%2�S�S�f، �IچE:�H4�&���O���u�lzC��9Y)�ɳgƂy��B�	�.���,D& Z@�*E?)<�B�Ƀ˾q��	�,2�>���H0f
zB�D[�#p�1C$z�)��[jR�C��4���*J9,p&/^:�!�dLT�d��CZND�qKP,V5aB!��9�p�v'�0/�>��V*�+:!�dR�>�J�A`�I�y�i����1~!���W��0�N;w^�i� Ch!�IO�����׊Zm�m`� �n!��(3j�-�;:]D�s  �!�䓍^�T��m��sN�\(��#,�!�d7���c��6�T��3�]w�!�d��`R����M�N�i)���PW!򄐐x�]�W�Ңx�$$��XbT!�ܒm���7���D0A��:g!��З)_~�����3:�b�AЂ�g!���*4GN`3�D�"E�\pKs"8M!��߸gz^���G�S��d��"Ov ���q���q��(�tHh�"O����% L�yH�c�j�܀e"O�1��M Y�,��P�̌�"O����L/ �1���J�$�d*O��eO�c�PA�]9iP^���'C�i�sj� >*���u*�r���'6p}��'ZF�0� ��L�d�>�Z	�'<\��.ˣg�6��m�X��ؒ��� ��Y�mܲ\9�������jp"O�ZVė�gN^<3����G�����"OT�y�����,���-Ǽs��v"Oz�;`��:H���,P�#��="OLY������P�	.۬�c"O�0�N�C���w�]�-cyYW"O�Xp��ε+O���$'K> ^h5�V"O���"�[�q��,:q�ŗP&E٦"O�2睘�>Xx��W26�,Q�"O
D %,�N\�Voȟ� ��"O� P2�XZ�����+\�b(�'"O`Ԑ�I�x���`J�
��d
�"O���n�/O>�q�<�\!e"O���у-b� ��[6w��K3"O��ZUcV�]:���P��"hh�*�"O�A:ǣR�A@�@�E6��"O
%��oM1?c��z���#�l8��"O�,���Q�^ř5Q0ݢ	JE"O�Ѣ�n:[�ҤpաV	,��`�"O����D�9���v�1"B��"O,1�B,ٹ]nn)��˔/6d��"O�z�,R��q��к"�f	�T"Ox\�sǒ�~��C��(�(�"O��w�ƪU^谰��%���B"Oxu����Lr��R�

t�*�B�"O��4.\���\���
:	�N���"O�4I#(����ĥC ^"�D"O�xCZ-���IՆ�jLr �"OX�����Y�4ܚ��^�vg���"Oބk��Y"vE!#Q�_]�l��"OJ�2�	A�b+�(v�n��#"OZ ɴg9u��"�� ����"OxQ�@�l�>s� N��@|��"Or�aa�^u��)�Ԑoʈ#0"O �е��//��Q3�9R^E@�"O�Q�D��6�bQ+��	6� �"O d2b�&1|�IA��>��a`�'��@���	l�֭��@W0��'M�#�лf:Ik�d�<(p�(C�'W4���ƃY�[W��Wt}��'�>��g_�#(�y��AR�����'�@ 2�h�a�|Φ���'��|�b���~�QY�hI#n��'��A*��Vd�B���Ε;�'_jE�d&ك]�
 ��Jx L1�'=�\)����F�I*Kz�F��'˖TC��M��œ�������'�4�ŬI�G�x�����c�`���&\� r�d�[�ސ��,W�~��ȓ<�����
[na�Lv�ӨQ��h��S���`'	~�\A���0$8�T��yz|�gh��$>�Yqրű�vņ�"Aр��q���Ё�ȓ#���R�b��?;�I`��r�Z��ȓT&��q`ɶ#-�xa��<-4.��ȓm��K(g��)��Ҽ
�	�ȓ�d��d�ϷR���ٴ*�ܝ��/�`��Ġ�� �J��b��n4�)�ȓFd*T�_��DЄ�͢^�� �ȓ3+\� �!B
��b�R$�z��ȓNg@�T̼);�����P�hD:ԅ�&���(��_ct�)�G�ZI���ȓ.�|���h�z�J�3���T4��q��!H�M�����/�����S�? �i �N��h��!�L�&���"O�����`��ܶeڔ�Q"O"��q�2d��M�o�BEE�"Oj�2d�;M"���H�D[^ h�"Ofػ�X8Ȝ;f�y\�4��"O��Ҕ��Qz*ĻD`'��*�"O*�y��%^oĴkЀ��hzj�"�"O��7
L�Mq�P L�fhZd�a"O qň[�m��z�/ū���°"O ��o[�$+*��.	�K�y�"OY3� )Zv\-�LF+N� �q"OB�S��M�1���2`Ԓnل���"O�]��O�ut\�(w�]�r��tQ"O֑��7�8�3�ʚ/x��;s"Of�	S�S�`p>�Ai�!ib���"O��Ò/�7K����	4��"O���%T��p5��fZ�g ����"O����C	����S���r�j��Q"O8�p��@�K�����ρ�D�(�0"Or|@�ɑ�g"�Sb�O�N��Ek1"O|e@�"Y/H��Dȯ�<��"O�
�.@�T���i�ݱJ�t0��"O�)��-Q|�hR�e@:-Q4��"O�(�.�;z?��8��V�X:�H�r"O���$됈����S6D%@u"O�5��)��G�l��d�'��c"O���b�ܝvQ��"$��
����yBO��9����ꀈ9h�I�/�y҉�&Ȯe��OCD�����h���y���&�>$`������@��yR����x8Wb�?y-.��dh�y҉N���B���n�Ɓ��;�yb텩	c �Bw���^����`��yB�D�HX��#ސ)[VHĢF*�y��GZ�"��F-�V�L�v/߸�y���a.@ 0bӆB�Ե���y2��s�T�Ң7���R�y�� j`Y3�.�6���C��W��yb��1hp�8#%�+�8���J���y�D���� đ�5ĬY�0���y��8s�:H�C���7ϴ�1���:�yr�K�{��;�%Y2t��D���yB��${��$���+A�5� ��y҃��&�F1�M%pzZi.��yb"W�wS���`Ѵ�����y�	H'략y�f�2!���`�L��y���<W@ahv#܌Y<��CG,��yr�Ty�t:�O�d�!�y�ʈ9W�\a�AI�0�F1� ��y�X�k�T� �J�whuf͎�y��ݴ(9��QQ�=�\�[�!F�ym)W]0���E䤽�A\��y"�7'��$ǬH�1"��QW�	*�y2��6ut�ؑi�4�`���K!�yRڃ/C|�v ���"+^�yR�в)��|��"L�9t�B2�T=�yb �l��#��w=E�$C���yr�C߈�A�"ʫZ���Ɂ��y2�ѐJP��ӍDQ��y	5�yR(P-��H��;8^֕�!�Ǌ�yR�$`V�	k �0,�"T
1�͵�y�ݨ���C�
�T����#�y���$�0�I��޽N���R��K�y���W�>�6ѩJ��Ћ6�=�y
� �qH��;sFH�%�� �RQk"O�Ŋ��S?g��i�w��-�04�"O���	_�@2�͔*���"O���.��ԁ͂��<P�"OLU3v��)�.؈��O9�"B�"O\ȷŮa�$q�g�9m��ҷ"O�(��(+|(r��/s�9��"OpH�&�/~��qz���T����P"O���ؔA�`�#Ӆ[�3�2�"O���7�V�+A��I6�&e]AA"O4��&nɑS����/AS\[�"OD�:�l � ]<i���M6oZ�6"O���o�g%���r ��a��3&"O��)U.�)�r�����GV0C�"O8Ac��"C����	4-���W"O��ь�o����D�9R�@�"O0q;C�M�'�P��M�� ��̑�"O5�T�>lQ�8�bT���"O��MY�C��8)�?B� �� "O Ń�[�B�t���$��4�"O�7JI8y� ��be&�T��t"OYQ��Z.���`���x�{@"O�q*V ���r��o&E� T"O"�!H8.���t�\�6{�z1"O�Y���?=�>����6^��8�"O�ةV��
1b�� L"t�D!�"Op%)����o���� ����S�"O�=8�M�n�����N��Sy6|�"O�u�k*v�3N��:PQ�"O.�)4l�`���i��g}��9"O�j�fס&�����+j�SW"O
|����@�܄
��U�[c Lu"O:�����N��<;�I�>~S:��#"O�E�G��_�:U"��O�����"O�A�́/5��9w
��~�=�"O*��ٻH"V��צOMeБ�6"O\`�qJ����Q��eҙMOƙ�S"O�h��ɞ� �C�v8�$j�"O�����(@�Qz��j>�I��"Oҍ��lW�
�b)�&d�
C�.$Hc"OE1��E�L�硋6~��"O��[�i�&Nv��b���l��1"O�I��d�z���p�zxc�"O�i�����v�pQ��;I�R"O؉��,�p˾�k'#P�o���"On9��M�&^�����H�>7r="O����(BP`4�&˧X�UcT"O��4��j�YFߚ�4"O\�ha��BoA�5�Z�y�l	�A�!�dN�vR~ȁ�@͓-�n��h��t#!�D�sL*�JGAȫ|������T�!�$���4X5�N4_z��&��"�!��I+��d�uK\4Bu�5��AԆq5�������M��OH����O��$iӨ�{�n�+@|M����%ibX����g������|f��{rx{Aчf�r�U��dlI�U'ɮg���i�nB����ɰ��N� v�čz�؆=D-z ��?1��I剀MCt#|����u ѧ�!LLXC�k"�Ҁ�a��ğ,&���ID�'��-�d&M<	�̴�u癮Em���{�,u�����O��oY�D�'ٛ�%݌O��8*� �]&i8�Q��~�Mљ6`�6�O�$�O��O�	}�JY�$+��L,!�*��i�J���%cڜ����p>y�a v۬�]5���E���Xi:١aP*��u���ևIP�(ư���E|���~��R� En.��AOD�s�ֈ�Q/�O���轢��[y��'��'��ia-B-:!��c,��!@��)�{"�'� H���x�z��#nҰ(q�m�!	��q%��`ش�*)O)Z��A?� ���RmZ�~JZ1�Q��=J������	g�i>��I�:�������#c�Ηh�p�$�M:+qj�ӶH8lO�u0�c�o�ԕ���(���]-E��qAQ*]�lRe��ɳ.(,�D�O6˛*U��.Up<�rG��y���ĩ<�����S'X9�Q�S6J�h�x�oZ�w��C���v ��A��l�A�t��6L>�7�lӐ}lZnyr�Ԗ�6��O�c?��CC�dx���>T�q+�M����I쟴���5�	쟰%>�x'(^�)Ŝ���a�,nu�epT�:���Vi\�`�:J�j����)VHu�yՆ�<d�)������O$��7�'��5�I�~�&F�������.�@��e�X5n=�O���<QB��5d�z���X�|�浓�'x?q��I��M��i��4b�����ƛ�jg�}`Rə�u�MS� �;b�v�'|�)����?Y��M�㝿w�p��%Z�y�0�Se-I6ykE�>�*���>�O��)@�J%j���l�Q���iC
��8$(������D�Yv�i>�#}�'�X�i6⋿x�|E�B$�$?����DO�Ov���Ԧ���9��>��BJ��a����ү[�!��i��ub�	m�'�j̋u�Fl�8p���U��\я{�N`��Ym�M���rڴ'��b�ǒ��h8�E�Ȝd?,���+	��ĳi���'tr�|�O�fI[)A�8S��Ԅ)��-��Pv���7*�j��P#c 	45@�G�1A�����k`ӈ��E�N�N�J�u�'�^����*_PS��S�^h����T�
�����O�lZ퟼�'��Z��n��
����PJ�.I0��ќZ��B�ɲ �ޝQ��J�<$R��T�T�ls�,K���d���'B�'��;J�`�� @�?�   �  S  �  f  j)  v4  d?  �J  V  �a  �k  t  {  >�  <�  �  ߙ  -�  p�  ��  ��  M�  ��   �  ^�  ��  *�  ��  �  H�  ��  P�     L � t � ' �/ ~5  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z�����W��K�L12$���SO�\1Yd�	�O�!�WR�H�Ī�.b�&hb1[��Q�|���T>�%		i�JI����z�`��6#1D��Sea�d]`b%�\th35D������?!�-Q�ė
?<��F.D�@3A�	5�Fy�B@WD&�H�!D�,s���CB>�rR�>dwA�*D�$0R�Ō*���B��30�)�-&D� c3�jFM �jp����('�ب�^��*�\�Xi��tU<Z "OlA�g`�$`&�@��I�kHH\C#�'ў�
Q�� P���]>�h���$D�\��.�h���p h�X�\�L-D������~`&A��K 1.V���5D�x�`ך_s��:��Yd8�4?ю��S7\�^5 A�ݯ�R=8�'��B�IP�&D���� �DU� �#$��B�I*1	@��G���J$E��LOO�JC�ɨp�\Dhfe�?`��鱺@�e��=O��i��b�x�Y�)[�ks$�ȓk��b#͔)rNQ��K�j>-����@�w�B�[*�� G<@�-�����DNA�R}�U�$���g\�܇��i��T}���.Ƞ��ĩ�C�(��C�	\?ы��?vԠ�F��K�#=���T?t���N�\Ry��:D��ۢ�b0t1��,�'b�tg8D����d�M{��CK,h�����5D�g�7Zr�#�o�!}�%3�B4D�pn\t���V͞؎i�sG0D��ڀK��/��r"�0�r%)��.D���u#�l<���`��MfNݲ�M-D�J���p���s�mX�1F�K7,D�PsC�Rj�����RLmXB%D�d�5mc�D��aiT�u:8}��#D�Da�H/6)bY�dݹV(Yxu�-D��Ԇۜ��e+���
Z�H�c+D��c[1N��A���5���R�j-D�xJ��S�u����@�b�``���,��h�4`Gf����B�f��C�Y�h �ȓ&4e�R�:�t�Bt���4!�ȓiW��
G��#�>L�s��)�z��ȓ3��Ց�B�	N)��ܞ.�4���o\\x��63X�p!Q��2����r��)9V	�4!(�E��
yI0��ȓN#�S ���(HG�ϭs�b�ȓM�@�y��/^��6"L�Q�ȓT��"��԰�h���֡�X��gX����H��O \�j��%g��ȓ.��0r��ݍ4�8�Q�<o]
@��I�L�Ӄ	"&^B���ǻ)�r���<�@,h"�L�\.t�%��6���+݆=s3��W���!DK҅��݄ȓ�z(��k���V��EU�j0���ȓ�R�Z��L�^��+��Q�k2(�g��~b��Y2���Mۉ\�����[��Ov�'	|�c)�*P�ӋA�1��Tr��,|]
g"O� t��v��,l��A�i�#�A�R_����)ҧ �`gc��Qq��a�.Jž�ȓT��1ٶKW Ĥ��@Ж3[^�%��z �'���W��-�:P�gK�.�p�'��Vhe����ȝ����9�bB�ɚC'B$XEi�3Q���R�( ����RO�tJ��BЅV�h�k�$G�n���BG(�<J��C;c��Ӳb[7L��09s*LO7/�I�QT�b�-��,r^ѳ'ɍ3?�*B�ɕ{�z�12LD�|��x9r�e�RC�I�f7�a��`� }�D�����B�I�5cZ����P9��S"S�84�"<�:��A�����Hy>���M�9#.�@�ȓC|��+t�/)<e@C��7hL�ȓ~��)��X9{���R��;'�<ф�J��,E�F)�prc��r���ȓ&e��[���88�£�8Mu�q�ȓ]o���1(�v�z���0rp���S��,�?W�Rqj��0)���ȓv�
�p��<@��x�t�������{Q����nU{��@�FF�����J���7 J%M��1)P ԂC�Fź]�� �5ݺ vNQ�a]�C�	(,�x�H �+��PC0!�)O�xC�I�$ޔreM�]J�s�OO�%�C�I��
��
�;.b��Q�����@B�	�Sh�H U��2d��vޟwu�C�ɐE������ ,B�2aA��j2xC䉏*hTŁw���x�ʴ�Z�}NC�	=<a��j�#9ZB [,W*�<C�I/odٚ&KиO��32j�>C��妰pb�S<(�6���'���e��&Pb���+ƾi�0ES���|m���Di6ʄD44$�[�oI0�^���>͌�*R���+�,�$%`��&v��Y�G�D���\�kڦĆȓ?8��(p�-^`<E�.��d��,��2B�ܻA������=��ȓq�*M30a B��r�
Ѭ��ȓ4ᐥ�$�G� ��u�s�x�\͇� xp� !�\��Ӆ�f����\6����?O����L��$�\�����I?e����$BXQc"O0�t��~�����L1}0��{�"Of�����x_y�3mυn(D���"O��ue� .��AQĂGT�c�"O�к%'��_�� (��N�;�>-)�"OT%���N=$��0f1=�Zغf"O�3�ɒ�}��%E��_��5"O ��g̓��V}X��ܖu|�1�v"O��h3�Ɨ$b(+����'U�)�"O���p��E�P0���s6�hA "O���1���!?@P��ͽ[���"OH�	c�$z���q��W�hXX� �"O�,�!FL��`@� ˭0@��"O���H��"�:�po��>:�""O&�h���Uc@��w/�uS�"O�9���N0�@V�r p�0�"O�K�b�g���9WE����	�"O��@��˜txs��u���:�"O*���e�j&ਣq�Ʌ:�xa�"O�X#`gE� & H�%�S���:�'�u�aL�ބ	������6D��2�gX�Fl�!�fG�5N��e)3D�� xk��+�:��Ç�'���d"Of%k�߃3s�l��On���"O�0;r��(A0E#�Í�5VΜ��"O��炍S��(� ��Er��J�"O�첗������*ݜA�Z-���'3��'���'b�'2�'�"�'=Ҹ���O�:�
9��pxF51��'V��'���'I2�'���'B�'X�)�w˗�c��] �Λ�c5��0B�'���'��'	��'���'}B�'���[���,8xT�,ݎjڌ�4�'R�'�B�'qb�'.r�':��'}��[ 
жO>^ԋ�6	��P#�'�2�'�B�'5R�'��'���'�0T��ˎ�uW��a�h]�0�4=���'���'���'b�',��'�"�'��\���l��Fj��JM��':2�'��'��'��'���'�]C@��'k�����^;P�����'9�'���'T��'H�'���'QlpZ�D���'���l1��'"�'�r�'+��'��'�b�'x�U�As}�IE���Z����'j�'ob�'��'k"�'�2�'d�ū� K;6\d�C�[�aNİ�e�'4��'���'!�' "�'D��':43׮�Q���jҋ�"dR����'�2�'�r�'jr�'���'Xr�'�8�[W�+&WV}c��C�H0��'���'-�'{��'���b�J���O4�I�;'� )��ܒW�L	geCy�'J�)�3?��i��M#Q$߼P�\�8T��4p%��۝'D�I	�M�R��>���`�䉈c���Lt�q�����
��?I�&��M��O��ӓ��I?�f�ޡ]�Ѐ!��_)�b�f/�ԟ�'��>ũ!��7��;ƯU+
n��s����D�<I����O��6=�QcT��� �z����:Lbpͺ�"�O��e��ק�OG|��i��$�8eђ��9@8�YWEL /��q���uUƢ=�'�?If%Y�0��&�;K��`Պ��<�-O�O��~��g��!GҢʂ��@�	�mS�2c�>���?��'��ɷi��(��K���#�k��9���?�ă>s$��|���O&����Z|����De�J�#W�'`�U�-O�˓�?E��'Ij����;�
}�)Ij~�9��'
����$��9�?�;Tb2h��� JM�`k�Cݺ=�����?���?�pe��MK�O��S$� -@.� �H��\�h5N�F@�
?# �OD�S�g̓Ħ]� �9q����������'C�ꓚ���O��?F� �nn�!B�����9Õ����OL��9���M�;v�|U�ȉb+R(N�H�l��@��U���D[�M�&�O@Y*J>)O�r�`� SF쁶���ļ�;���O��$�Oz���O�ɯ<a X�\���t��Qjt�ܻ<f�X���D������/�M+��>����?���;q(�!1c:�ȣ��]$J�j��W��M��Ot�X�ʀ��(���4(H����ϑ���"�l��-�$8�O��ꅍ݈P̶)S!aR�+��Ai�<���Ss�)ڷ�i��'7��3��DD�X�,0�P!�!VM�	ԟ �i>ug������uGʜ�4&,`��ေt0X�A�����[�'<'�ؗ'���'���'�9S�+?0�.p�&V��r	���'�"[�D;�O ���O�D�|�!�!+�x��C:��Q�`x~"�>Q��?aH>�O���c���
��<����621|�:�-�.&� �B�i$���|*u���t%�H�̌7c��%�CȒ��3&�ןD�I۟,�	�b>�'#�7���I?�e�Ч�wL ��>.��D�O��d�����?Y0Q�����iC��yu��+T�PX����6˞���ݟtj�cæ��'w^M)*�?Ť�܌YÁ�
x�^������t1O ��?���?����?����I�Jtԝ����=��Uq੍�/�y�'��'a���'M�6=��)�YY��1�
�iu�Iic��O^�:���ʍ:�6�p�@�Ư��0�p�v&T�^$pUh��m���c��mc�E��ty�O_�Q�z�{�(ȣXw��ht`;_7��'���'Y�	���d�O���g>�!��X&c�2���xU3��+�	)����O���)�DȫP�qz��0�Z�{�[�D��ɣN��ٰ�����|R����ɻ��u��dC^�Q���~#� ����	֟���r�O�Ҏ�z�J�����8ت]}�""�>����?iV�i(�O󎔽{��)1̂�E�0�$�7���O����Ov����w��;��� vG�?���`��2��pH��� �h�	Sy"�'&��'QB�'��`��B�vK�$�wK�t4 �S��	�OV��On��(�)�O���&�0Ӏ��ܵ4�Y����k}�'��|���J߿<H������'="*�����d,`^P�"���OZʓ^��a`�M� /g�
ņ�:I~���?����?���|r,OhI�'�2BD�3H�R�р�\������!£f���p �O.���O�-�	���1\ǜ	A�*G�G�h���yӔ�y�I@wK�?�$?��=� ����%$t�zP�U	L�e2O��d�O����Op���O��?��A��B�vi��!�~��}hB�ڟ|������O��>�M�M>���]�8H܁���,=�9��<�䓜?��|z0��$�M��O.({U�ŷ,À�J4!�w*��� �E��rx��'��';�I���ڟ���62Ƹ#��]�)54�B`jC�B-�}�I��4�'\v��?A��?9+�Np�rϽu��2�P�2��iR;O���k}B�'g�|ʟ�8�B��j@L�2�	�HD�S��ԦyZQ"k�`���T��K?qH>9�$�PqpD��U� ��p�B��?���?����?�|b,O��m��X����+g&aH0��d�F�	���	�M;�B!�>1�s��	���{���0G�-8LP���?���M#�O���ea���P���34�*A(A�8-�e�`�,�'8��'���'y��'r哶2=n��ˡ=L���	}vҭ۪O�d�OR�D:�)�O�oz�c�!�:n$S�]�j���S�П���r�)�,�n�<I�	Q�7�0��f�6�����J�<i3MHih�$^.����d�Od�d'(�Za��k�K�hPacd�/j ����O����O�˓C&��ʟ|��ݟ@��+ L��XF��@���U�8`�	����B��
���ȄX.|���è	uC��\�-��@�&�Mp��4āA?q�,�ʐ&ƜX��`��Y�S�8�K��?	���?���h����� ,�h��R7R��
���eB�Ą@}b�'&BBb�N��]G�>u�4�-
]����3J���I�����̟�hbA�Ԧ��'3p���R�?��4&δ�;"&�8&\���H�6b�']�i>���͟��	ڟ(�	�xW>����;w:B ql�Ґ�'ߠ듡?9��?iO~*�������I#S44h%�߫j��-9�[���I��t'�b>�&��9 ������䂀+�)Ov�m�`~��� �>9�������;V�\*�f��G�p��L�-%TN���Op���Ob�4��ʓ7"�	���ϨLh�Ɉ�@��1�V�h�8�ٴ��'�N��?a��?��:B����Մ��(��)C�|�4��D�!�����'f疓���N_�����X� �>%�B	�"p�d�O����O��$�O���3�#sB�\0!AաQǊ�2�+�[O�<�	ğ,��%��4�"���M&�d�TB��x��(0dQ�u��0:ECFt�I�0�i>iac˦��'�,EP�IN�~+�@�����9[�i ��¼����&Y)�'��i>��	���I?�( ۓ#N\ЈeX֮Št�	��4�'.v��?Y��?�(��kj۞3�.`bn�0u��\r����H�O��$�O��O�
��E�LL�36~�*�Q�A�zu��\��Z�ls~�O�\����%.5��*�?X@`��6 S^j6����?9���?��Ş��D�Ʀ�3t���/@���L���؁�g����ܟl�ٴ��'{F��?i�&�Rʀ5�WA�|�>��˔�?i��ed�޴����2w��Z������Y�0���(k&x=�5�ˈ�y�_���I|�I�\�I۟�O!����K	�G�"��C.M��y��>���?�����<A��y�o�9j�Y0&	# ~���5&P�RX����D���6�j�pàS(Q�앛c��
�r�h�*s���ʞ�8�)�M��{yr�'��Y�	t���I�<W	 }�p� R�'���'^�	����O���O����e����y� �%Zp���*�I���d�O��D=�d�l$�����D�N�B�鞿Q=��%���".^7��-'?I�R�'��	���X�\��1ᇳ>�ƱKq��N����ڟ���ퟜ�	b�O���G?U+TA ���f��=�煘�-&2��>����?Y��i�O�#Kf�L�/.?�h��QT��Or��O����~�*�Ӻ��7��d&�\�r�+qƘ'[����-�B@�O�˓�?y���?���?��R�P�����e׺5�3�[� ��/O���'��'���I�=b���P,�+n��b�G_�4��'	��'<ɧ�Op���,^2'��3��#dQ� ��q�֋�<!���J���Iu�eyr*W?:��2��'"m��a��'PR�'d�O��	���d�O0���P�0��P%��	9L�O�5m�h��r\����ܕ'>��/v �1�/:�)5�!L��р��i��� F�0� ��Od,$?���#:�����P�-:��cb�I͟,�I̟(�Iן���H��dNX0k�gKQV���a"aurpc��?Q��$�i>����M3I>!�n��~����a�
g��I�7���?I��|����.�M��OJ��f��"��"��ՋcJp�S�Z�r�.9�'��'���韬�	�� �I�I�Ķ6�jh�ɣ��[:}s
`����ԗ'؈��?���?y/�
�{� G	b8QBa,>)�hӕ��*�O����O`�O�ӛ��T��ˈ�|,�� �'!���0iO�|R���W�<?ͧ3����C9��t> �WĜ:8\���  �	�����?���?�S�'��d�Ҧ�	7V�eN��Q�-wܒ���)c�D��ɟh�ߴ��'����?���P�j���J�	o�m+����?���q�`i��4����*����mk+O� l!�s��!`1^�����g^��9O"��?���?Y���?������<���P!�}���`��(�xh�'<�I��0$?i�I��Mϻm8Z�Z�o�m��	A��Y�b3�����?�N>�|ʷ��M��'�X�ZQ@�5�(��DȄf��q2�'��Zc˂��dhƙ|"[�t�I��l�T" 	���ڂ4��Q+f���h�I����y���>����?��ф�qį�V��R�(�<�@A����>q���?J>Auj^2�6�9!���7�P�R�K~bBZI@�I����OB��	n��+P0C' bfͺ:rN�9�-̉j�2�':b�'���S���c��i���6Dͷv" ��6a������O����O��mZ]�Ӽ�iә��"���-��XFh��<���?��8:����4��D�-:֘z���u��B4uT���5��M{dƐ5����4�����O����OR��n���f �2.��>	���D2����I��&?�	�q���b҈�'{���*�a�.H����O|���Ov�O1�Ԥ���a$��c�Ӝ]�J��2J��*%�Hv���
�`ԼUP2�Zr�}y��?��`�y`�;d�C4���'q��'��O�I����O�,z�lV����!p� ,����M����Ħi�?�P�����杚^��1�4e�%7�T�9��P�E�N=�B�Zަ��'s�;���?eY�����w"�b�@�3��Qi5!�9����'g�'\b�'K��'��V���'�"�xY�O��-���p�	ҟ9�OV˓1O���|�0 �ưX6(� � �B��Ø'+BU����U���'��������^
K�D|���M=����'���$���'!��'��'s2,z���\e�s�T�(�I�'�BS� ­OZ���Oj�D�|B6�Ј;��j��$+qp��V�X~�,�>���?�H>�O`����O�ډ�cX�B�XQ"&έpsl�ˇ�*��4����Q��O�I��˻���p�7�rH�I�O��D�O����O1��ʓX���@�P0��#J�4}4�A����yB�'3eq� ��ѬOr���'�lUJ�\]���S�+#(���OT��c�m�,�Ӻ��ޓ��S�<Y�O:˞}cрˑhb����%O�<�+O����Ot��O����O�˧k�� ��
>�� 	pN	��p0PU���I��8�IM����������`GL53ۈ�ׁ�0_�����?1����S��T��¦�����YH��W*�"W.<%�FEC7�y��V�z��!������4���$�x���ՈM1@�`ʄ�
6w�h��OR�$�O"ʓd��IKy��'-0�]8߸��ѯ�W4n���|b�'%L��?����H�ʥ� �B@��h�j�� �'��\A���NS4 ����D�@�(��'��A8u�P-:Y��Q�_�a�I�����͟0��p�O��#G�$T�y���>�ԅi#d؛t3b&�>9��?���ie�O�E3;�6�����.��hE�9_��d�O����O:ݓ��b�v�3�DifN��� ��+�t�X"�4	� A��\2�䓞�4�`���O:���O���j����j� �m��F��˓K~�	Ɵ,��ҟ�&?%��3֢��� G>��g��\e���OX��O`�O1�U��� Q`n��ED?8��18�M�/Ȳ7m2?�� �,���M�IWyҬЮ*�:�:���C=<�(��΢n�r�'8��'M�O��I����O�����"(��@��=QGt8"��O�in�@��u��	�h�	П��KN�C~�Щ@��y�V,�f�ٷ1ъ�mZc~��g�n��]ܧ�����3^dd5����������<����?���?��?y��d&��>���&Y�s�=��Ob"�'a2�>�'�?Q��iB�'&~��q�"+mrh� h �]y�Ĳ�y�'��Iq�BLmy~r�Gm�*�a7g��+�keh��#&^�dq�|rV���������ʟ��Р�q�:A��.T5E\wc�Ο��Ipyb��>���?�����F�&~�L:��L?x� <sD@�|O����D�Oj��+��?iZ 
�q��xR�[8���g�����A)U�'O�����$������|����F�8YǍ�
i�����I\s�'���'����[�l�ܴ��*��a�0���n3�f]�<���?	&�i��'m�>����d�q��vYj1�԰����?A��ߢ�M��O�N ��x�I���$V��T��==a�Z��4)��'@�����	��d�	Ο��	\�T���}sl��Ւm.Θ�2��-Db�����O䒟X�d����/#�g�ƞJ�I����nh�x��ȟ�%�b>M��A��ΓrDX4IG�^�*�X}�2F��X͓udX�"2h�O�h�H>	*O ���O������3�RYP��%�.���O,���OL�d�<9�Z����̟T��/#*�K!��*$��A��iڝ|���?��^����ʟH$�x�G�O�Y'��4.[�Cw,a��OTdʕ-�V��E��"�)F��?����O:����m�*�j.]�^�6 c/�O��$�ON���O��}��^� �cZ�/�����"R�����	ȟ��	�M���w����NV�-��'ڳ:0BpC�'�b�'p���j�v��ĉ�����4�>� \��D�K���vh�Yn4�A!��<ͧ�?)��?a���?�'��R��{�Ġy�(p����ċx}��'���'l�O�d��)}��Kƛ; ��c��0`D��?����Ê;p�XR̕��ܱ���-3A*̨f�\���?w��(�`�'7p'�,�'�p��΂�)�.m�#P�%:�� u�'�b�'Z���O��	�����O�5�͇�=�xX ��5#��|��O*�mZN��n�	۟�����8����ME��b�L�hLfEȠ�A�t��nZd~!	��lD���w�Ĥ)�	j�)�Cգ#	�(��'m��'t2�'�r�'��>)�➓�N�G+	�f?�qj�<Q��<�i>�����M�K>i�넔{u���bʪ���GK���䓲?���|b�W�M��O뮏�sԤ��/Ҿ��Dz��ʲ7Dވ�g��O6�I>�/Ob���O��D�O.1�P�XT�:U�"&*,�,5�v��O����<95S���'uBY>� ��F��rx�GG�/���g-:?�5Q������$��'�Ҍɣ@W�#�Px��H.O��<��(�����KDK~�O!hI�	���'��ݣb�?a��A�p^8N&|�v�'xR�'����OD�� �M[`S>]���bꎉӖ<���<����?q �i��O\L�'+�m�3h�+��ZnЬ�����'��g�i*�I�J�cq�I��GZ�(��~�F��ƅ��K��<���?)��?Q���?,���� �
�~?�!�g�4Fʈ9�O�V}�'y��'��OxRdn���!�4��!
� o�q�(֯T���D;�)��06Lao��<q��l�ܓaA�<E��G��<���=��Q8����d�Ot���&��p�LVK��ェ�\����O�D�O��r�	����	؟$!ҫte�BT��c��9�
@-}E�OE�'!R�'��'QX��0%�6T`�Lإ�S�!$��K�O�4��_�Xe�py��,�?)��O�X�������ܼq�,��en�O��d�OF���O|�}���'Cr�)��Z�(zTL,U����Z���⟀���M�M>Y�Ӽ��K�aw$(���!Q��Y���<��?���r2�1Pݴ����R������Aa�K'W��0c��:S�ȗ���䓺��O �d�O����O<��A����WK�� XS�/Ԓe��ʓ)0���`�����%?e�I5s���xF�72f���/];~PDջ�O<���OʓO1�ִ����V̫�@!�`y(`M˱P��7�+?��a��(�D��J�IUyr����} ��u_bD	�	�+xJ��'�"�'��O��ɐ����O�M��ݼjC�!�$��CT�L
���O��oZr��p��	�X�I�ɰ�Ӣ{����B��cK�l��	S�p|�-l�a~��*Lc0<�E�'���E�fN^94� >
EP�0b�<a���?9���?����?���$d�{�oЅ�^��ah�e[d}*O&�d n}�O.�cr��O�=aU���h@�Y\\��!�+̮z��'������<e�6�0?9�S!*1f��a-͇!��)Q�GR�M�<M���O�|J>�*O�I�O��d�O���M��@�ҟ5;�P	�O$�Ļ<a�S�X����|����cƇ6��"�ӱ>�0@�����Dc}B�'��O�3���$M׌;�	B�]/e}�t1��؜v���Ry�Oxb��I�C�'� P󂓼U���
ˉ\p$I�'y��'�b�O��	
�M��l� A�"�� B^@�Vurs�E�<	��?Y��ie�Om�'SB�QGyD���F�7M@�4c1�' 8y��ip�	Q\��Y��I?Z��m�5Q�_
x
%��G�<Q���?����?����?�-�h�� ��.��0r/ʅq}�(�c�Pb}��'Pr�'���y�es����A�b}ӄ�P�Qh:5�P�$�O�O1�v}�Kl��扁qs���t�0 �m����)W�物J-~s�'�θ&��'���1���	�Hϵ��ta`JPY������w}�U�(�ɯ8���C`�_�lh¯̑o^���?9�\������ $����%�5Qo�h0l�`6	T5?9� ӌG���˖��O����?�Ǥ<fQ@��-A2K�4�BSeĔ�?����?Q��?y��)�On�["�*|���Tk��iWd�OY�'���'�7�0�i�q��e� z7,����!��y)gh����ڟ��I\��<n~~�j�;pQ����������� 0B0[��:��u�a�|�[����������	���"$�c9v�zGOV�;�X��c�y(�>A��?!�����<�dőE;<��b��B�B���#�YG�I���?�|:Sl[CҰ3#�- ]�D�G�<���2����$&�Z�c��4ΒO\ʓ&v��p��_�,���+��xJ���?A��?1��|B.O�'I�e����Ӱ#� ;P�d]�X"	�b��J�O"�$�<�`��FͺtZ%�O�^`�!�o	�/�����4���ľ>( ���',�F��8��τ4����@\�Z5����*P���O����O����Od�$"�S�{�l�h"�˶{H�Q�ݕ���ɟ\����$�<�g�iW�':��1���A�Aq�.�5�\՚�|��'-�O��9P�i}�	� =�� R8�5����(C��&����#�? ���<�'�?a��?T�@�3��<p�D4g7P}��C,�?����@}B�'�R�'��ӍW���J�f�fy���U�]�v�|��I��\�?�O�h|��BOgN81YA�윳��F�|v��Ē
��i>m��'N*&�T{@��?r���$A�;��Hc�P��|�	�����b>��'�b6�K&�EB �?LA��e�Lm�<Q�i��OTA�'�r�Y=x�x�v��4p�f�y�&��C��'�<A�i����&��M{`�Or�&��DBΔc�
삢��'��<�,O��$�O��d�O.�d�O6�'>w:V�E�&�� �V�lP"�IR}r�'=B�'~��y�Ga��nܭ~��aH�*l�*Ex��Y*TqF��OF�O1��UX�r��ɏ\^�(*���e[L�"v��an��	�'��I��'}0-$�Е'
�'�P��$�{�R�"5���{�>T���'}r�'��X�0	�O>��O"�$A��~<ӶB��6�䭔O��z�O~�D�O&�O ��w��YZ<��(՘o8�����x���<O��pq�'3�ӿO�'S��JQđf�ĨH#oDh�D������ٟ�	�DG�$�'�*0Ҳ U<��3`�6&z����'=.��?���S���4���(Go�)OodB���b�DR�1OF�D�O(�䈥p`6� ?�D��4�����M�D�8��Y�pl�К@ �4J�8�%�ؖ'j2�'@��'�R�'�@���B�T�Y:��)�l��_�T�O���O��=�9OI �,1��ʦ��m���@}"�'�2�|���MM1V�3�#�)�-����a�:4s�i�dʓ���!���$�@�'���PK���X�%�Q�<pRB�'���'7����Z�p�O&�DZ���I�`�L$�*����o4�D���?']�T���X��'e�4��TH�0�
���5l��Y�CԦU�'԰�B��	�?-�}Z��S��Ab�H�Dt
��OC�IpΓ�?���?���?)����OnDAzTd:?����
�	up�K�V�������4�����٦�$����1~L���[�x��cq`Jj�I����i>��W�AӦ��'�j4;��P-�łD�cQT4@7��8!�l�I�Y-�'��i>��i�MS��`ʜq3 �VcF�b��5Im�����?�/OFM�'N��'^RY>�j"�I�5lpzpꗬz�,Q �e�H�ɤ��d�O�����K$�Q�!(n�ha䆋d�p�!W�D��@��C���'��4+��!��|�JQ��y�GM�W�*�K���e���'t��'E��4X�hbٴtf>�s6!A�K�vEZ1/�6�����?���v���|}��'*���#
�v�p�%K�v��M���'8�A@>>�摟֝�r��Ӝv�割>�D���o�QC��R~
�	@yR�'���'��'��[>�hR	i�|���5|y	gA���$�O��D�Op���������1o�<��� �)2H�u�2�v��ٟ�&�b>ᑵ��Ӧ�ϓ4��(  �	?�"�Y)z� �  ڜx��O��䓄�4����]�Xr$��%��-�zy(p��1eמ��O����O,˓@��I�T���|)t�-���kV��-iC�W��5|��ş<�IX����(�L"� ��O4RSF�E
\A��I�Y��@�|:���O�@���Jq�j	R��1�R�I�.���2�L�O4���O<���Or�}z�� ��c�N�wd��6��&&�j��xg�Ipy&{����:`br�� K_'	�v��v����I���	˟�yO��)�'.��p��?��a�ܤJ��EO�R�JU[��I�l7�'��i>��I�x��ğ�I�>���$�~�i���(���'e���?!���?�J~Γi�\�#���v���lު!$=��^�4���%�b>�O߁$S�p�׾<�,y)�e�I��>?�R&���<�d
=����	!|�b��sm^�*yv�i�ҝy���OH�d�O��4���!]�	ҟ�fl�b�����>db1xD,@Ο<�޴��'/���?a-O�R����ar�嗿	��&�Ϗx7M!?q ���p���iD>����V���ٳ�ED[�t�m�!�y2�'�r�'��'r�IL�v�!�V�; ^Q�E�����Ot��j}"V�X��4��B�l�Bg��>.1�<�u�ŝuF��	L>����?�'�� ��4���P(3�`�DB��3ڬ�Hu�^���D'B&�?i��:��<�'�?���?	G��;&�P�3��)��[&V��?Y���D�W}��'���'��1�D�r��,Zq<�C�	[	���I��Iٟ���b�)jt��Z���aJ��`",�:��RF��7MSk�V���ӮrC�@�6��-*�Q�Q���L��\�e)��|�ȕa��6�1���*G�ʹ`�M�J5�X�}q4���+� �̑	d�K����E�?l�b�*ƭ��b��ׂS)t�����-.�K�]H�Ξ
J��Y*r�_�0��=��)�������R�����!�*�[ ��"O�H�����; $a�+��3L`�S���f�06��9:���4G��L*ŬE�k����3I,s5lې�ƩH�Tڷ�X�4����B4 Ű$s	ιg�fm�p@]���S샋T����
&C�:�@B��*i?���>,O��D(�$�O����3)�RM�V���D��C��Jx�*�O���v7O����O��$5�ɤ?� 4�2�DH�y�1��Oh��H��iCR�'��|B�'�8`Zc/L1a�"_fPh����~H�X�-k�����4�	���'9����4a��W�~��"�(�3n���f���M������?��cNT�a�{��J� �$��� 6p�8��M���?��+��<A�����OB��O9��F��iSk�!����Ң�G�����ɔk�r��?�O���N�-Ee���&�X� ��4f�<T͓�?����?A���?�����ٸ9M�����P�|stI�%4���n���	��nm�?�O%�0*�4cHʂ"ۄ:�$<@#.��l�ϟL�ش�?����?���m�	Dy�CҿR<���	�g��c��ņ�F6�����D�OzH�'��ē+T�^��^��68��W
6��O���O��A}�W�(�	}?!vN
�aP�5�B!ά3�"����FX�x������V�x�Γ�?����?��dH ��h8� "�h�&�M�6�'G�>�/O���5���<�{��X|�T]i2 ��M\0��R��7J�ҟ�u��|�	؟|��f��H!p�v�у-[OyR���_!���ly��'�'k��'@�����2
 ��ӷ�C1q���kCh4�y�-A��y2�'��'!�Ol���E������j���V(E�:��7m�<	��䓗?��7-r���'3H5�"�L�E��Z���lk�L�	���	��'���Op��My�`$�,��^�ؤ������	D�	ß��	���=���[��(W�_/%��������Iٟ�L{������	�O����Okǧ��%���:4h8�%�A�cF�'t�	�L��L�s���!�� ��
��zrT�S�	~6��_���Oh�oZ˟��I���	7����3jq��qk�'6�Z�H",,�V]���I���aI|z+�NM��iμ��`n�`s2%�!m�k�D}��'��R����KyʟHH0fY(��Z�FQ<iG�` �W}��%�O󩎃��ɾ�𥱢�N��=��]���"ٴ�?����?�����?a�OH�����S��Y�w� &1��qk�_[�'�"��z����?�Ӻ{����1�r�R��:D3"�[�IĦ1�I��|�'� �'��'�	�GǛ;��A�cһ>"t�Ƨ%��ҹ5��$�����S_?��C@�.!�h�ӗ6Hz�!�
��'�2�'�Od�Ģ���2	�*`h�4;��ľ o<E�Fnt��|���.��	�X�i>��'���r�P�
�F��Z�XM��ݴ�?����'W2^�P	�&dӐ�3�`�/k�Nq�)I��n@+����<����?y��M��O�8�'�?!� �b�Ȭkc	0�%+��Zm�V�'��'��i>9�	B�	^��^Ţ��Z�T���Xw"GvW���'b�ʇn��E���'����56�M�[B��P��(=>�m��ē�?�/O� �u�i�U3Qb� �2!h��(�n�8�FxӶ�[�;O ��
������$�	����O��`F@T�ZY��*�d�i��`�7�i�����I���'��� �EÛ��iOt�2�.�!T0��`�n���D�O����OF���O�S�Tc��X��lޑ"�y1$�&Q�0�p�Fx�OR�ʛ'��(�A$P@#�
B�6d�!Be�"tn7��OZ���O(��m�)��'��IKhH�/'��X��5t��,�ݴ�?!K>)����Γ�?I��?���_����A�d�0��t�s�7S����'���=�?-�'��� Q2�!v�-vg̫o��'�R'�y��'cB�'��'')�I�b.A�~)��YA'���2�n��ē�?���������dj7��?2ZuA5��@.�� ��i�b���y"�'=R�'H�O���S��\��$�+6~�� �A�^�듧?�������4���Ē6���"�طx_��J�;FWN��0O��d�O��$o���I�O���C%��T����hY�9���æ��I[yR�'l�'-Dq8�O�i����C��Ѕ�w	T!$!��4�?9�� �|͓�?1rY?]�	ğD��/JE�P2�.B̙Y��T�x����O*���O8��&N����O�ʓ������e���/ �>L�c��	�M+dM��<9�x��'���'�Bm�>��]:��qD�%T��"� �d��o��l��}��IZ�Ij����M���L�'7؍ �ж[�hĢ֊Z��y���M���?���?Y7R�Д'_r1�t@�.]�0��!��2�R�}��	�<O0���<!(�ƹ�v<�b�D��J��Xs�ɴZ?���E�¥0$o�ԟ��џ���=��ĩ<���~�̖b�����=r.�M�u���Mk���6��$� ���O����O���h?2H<��TwG1C֏����ߟ���O(ʓ�?Y+O*��ƐDZ�-�6����獤(����_��D�}�����H�	ȟ<�	�?�i݉��gXz�"��aCͿ:�����{��'>�	P�'?b�'	�J��V"�JS"�5T��H����o����'����'���'<2��$�>y���)���o��!�,|�4��?�/O6��O:�d�����1Jڢ\�fI�Ch���ٻcE��X��'W�'7��f�m�O�n��?�1��Т�H�쮁��c����l�ʟĖ'���'+�/�)ߘ�M+`Hϱz�ʗ^#�=��/U�H�7��O����m�D�O$�O���'���8� V��$LbG�TSiM���Qf\���ʟ��	���	sy��'���L�/p��0H#2�ظ脖ś���y��'�7-�O���Oz�`}Zw�SD�Nd}{V�C�kV^���4�?���~��������u(��$U�g��R��Xc:$�ed�$�M#��B�6�'A2�'$r,�>I*O�<�(�!����.V*�!�B��Ѧ�X�%p��	yy"Q>�92�z>����C��lanӚa�l����e�V�ٴ�?��?��&!��Zy2�'_�d�3t���Ȅ1g���Ӷ�+_���y���yr����t�'���'��*A�fz*�A��Ǘ�>u0��n�"�D�O&��'v��ޟ �'wZc��l ��a�0���	p�D�@�O,�&2O�}��%�OD��Ov������B �ν1�sW�do��d�i�f����O�˓�?I��?�/��}�~qdT�&t��kdfE2"�Γ�����?���?yO~3�����-��EDN�a�#�)h*��V�x��'C�'���'�Zՠ��'߾���2D�5p���e:��*`L��y�'���'8*��4�O9���=y����Ǐ�-rݸr���pP�7m�OړO��D�O�`�2OH�'<���_��v�y�!�Sֈ��4�?��LP�͓�?YV?e�	ş��1cLL{���2�܍��\�`��N<���?��b��?YN>A�Om�,�GM̫t�5�R�W���`۴zVt��?źiB�'���'X^�U�Ri�q�J�YQ�� �Q!Sr��m�X���
�x�Iu�)Bq��Ӧm{����	��0��Cx����z���WզI�Iޟ$������}��_�L��S�j���Ē{�B7m�'&Ph��#�$�|2g�R�<I��i&�͑��+5Q�I�AD؜#�as�i���'=r�'��Op���O
��O]昳�? �]բ�=o�7m+��ژI��D�	��O���O���aO�*6S�1��.N^Ԙ$�͝���I��$�K<���?�L>��*� j�D5|D����4�&��'�؈82�'`X��'r��'�~R�-&]Hu���2�̆Ҧ8J<	���?�H>��?����� Paǋ�\b�囕IT9P�Щ��j�B�ϓ�?a����OH��ST��Asr�S�9����S�P,M���?)��䓡?!�y���x�Z�X�b#�
6��A� Kk��¦�Ҽ�y��'���'T���h�OU��p��a��^�I��dx��,��6-�O>�OH��O����:O�'D=��(��^��3.�&���4�?Q�I�8xΓ�?9W_?M�	ʟL��{�m	`�S0����;v�<�!L<����?�g�H�<N>��O�X{��ÔIҡg�D�i�t���4pb�ϓ�?��i���'W��'Ϧ��0Y�˜<h�^%+���RE^)o����	�ut�e��j�k�����M��A��P唄�U�Ʀ���*�M���?1���?�x�O<F�0��7�ƕP̚�E#$�[���>�������#E�yr�'�����
=Z��&��(&���jk�����O����O�`�'=�	��,��r�:V�U>(
L�1����9m�ϟ��'{����'Ƭ�P�O��'��#�%ReԈ*��ŇJ��x�'	���6��O���_}Y�p��Oy��5ffS����@� .��������<�D0Og,�D�O��$�OH�9O�", ��(u�Fm�P%ߣ6{���>	/O���<���?i��2ۤ��w��m1Hْ�� �yۨ6���<)�lK��?Q���?�����)�T��'6�li�+,J��AM�eWNxm�SyB�'{��ӟ��I�D��Bk� ْt%LAR���9M,�#LT��I�0��ҟ�3O|z�Y?��It�9�Bl�<[�����CZ�ՙݴ�?�,O����O\��ٸSS�Į|n�Iʡ�A�0_�P������-g|6��Of�D�5o����OB��O2��'>�������xr�n�lAp�f�Q����?���?�C�J�<*��d�?�3ƒ$b�Ɛ��V�n����v�>�i�3O2��ܦI����I�����O��wJ��� �&%�E��&F
8���'���Ԫ�y��~�������y��΀�0��h�"��`���󲇊�?��?)���?y��?�*O��ER�H�'�]8y�IThZ�=R�\K�O<4p��i>鲣�e�p�ɲ~ǌ�`gI��RYfɳs����}�ٴ�?���?���37�'���'w��[p�J�C��q�ԁs@{3�� yT�o���ڟ���-8���EB͝3_����Y�(y[�4�?��P�'�b�'ɧ5֤
�qeb����Z�$���� �%��'�ȽÝ'���'R"�~*e�V:q�x��A�;�D� ��E֦9QO<9���?�J>1��?�-Y2{�P� �����;]I��Γ.�\0Γ�?���?M~��4����5��d�7�4"�d��`Y�P���\%�T���DJĄ�>Iö��)9UD'K��1��O۹Dl,M��?���?�3���'�?���?Ѷ�A�d@���tD�@�)�%-��ga���'��'��Z��ɂ�6�DO�V��xU��U�ez��̰,V�&�'�B%^�yb�'E.ꧪ?Y��?�E��&qK�LQ#!8e�	sЉ�KO�6^�,�'�4|�͟�I�?7�E�G	"�#���V�4<�d)�9�Ǟ;���'���'t�	���������U�d�STh�.R��Y4���M�����DVB��S�f��6M�}�t�3V��#}QF�2���*���' l6-�ON�D�O��_M�	��� D�$蔤8.ƌ���|O�p��i�����?��5fj�p��*A(ց�6MF�!���
2
xV��ٴ�?����?A�
;�O��䠟�C07e�T�8�1~O�m�VK%�	96�h�	�;#j�۟(�	��HC�`ܩl���H-��F�]Rt�+�M#��?��xb�'7�|Zc��D�f�B"S�Y�i¶��0�O��B?OH�c:O"���O�D;�t�V8l%9Tj^SM�J���M#��d�On�O$�D�O�d#&O�pu𨂳�q+�<��"���P�GT�$�OB���O��ɡ|*��5����rK�r�MZrѺS�Tq�i^R�'*r�|B�'+��/H�6MU/�|�����?|R�	��D�>Z��Γ�?���?Q��!�~Z�-��<�ա�
���i�Ԡ@i��Jֹi�R�',�	ry"f ���Y�8k�� �`Z��p�b��8Ґ2�Hg�����O�q��.�O����O��d�<q��g��dÌ�s���81��_Z��aƒxb�'��	�d�
"<�;^�(��AE=h� ٻ�Ą�R�\9���̆c���v���a]tX�UK�Qږ�X��_4{�py�Ɓ�F�,�pd�ˈ_5�`�AD�bt��oI���%0L�A�A̕K�n�p�AΔk]B 1�A�N,��Ym]-����8��s�W4R�����G�Y����#z��=�ڲ5E\�1čN3�v�wJ�&q��]�E�u�0��QD�(t`O)���EcңM��}�Q�F�T+�$R��-A^�z�kܪi4d��cH'㨭��a6a�s�ፘ�f�q0��;X*\!��S�C��I�B�r����.}=�v�'2�'���P����$��@���v���eK"a ށ#��#�h��bj�+~&��ư?�=�� �^�Rq)�ƫ>�y��Q�<hB�
f޶<�Ŋ%��Q�g�'f:8�׌G8��tc�7�����';����?y����<!ң�{��H�M��]�g'^�<!�m��<Q8�c�����9!��ۥM#���'��^�G��pm�D�� A�EĚ~���Qc2?���	ݟ<��Yy"�'d�2�t$��I`\��@\�	N�WH�<�,1#1cclr8<O������sʕPp.@#:f�h��ͅ@ٌj�Vr���� 0<O� j�'��i�bktأ�J.3���b!4�ў�F��@.��sĂz �!cD��y��.aD\�Á�*|���,ј�y�+�>y.O
ِKWt}�'��9d���a�@�FԉiRi�.���۟���������S��P���2'��|�RM�m��{aI�Y&��S7�P�'�С�ِ.�r�*%��~��JRe3o7�8��]�:�@�<��ݟ���'�:)� ��6in���S�d����?���ג%	�p0G.U"�p��@��rI<Y4L�.)�́��!p���h��<��J�}��ǟ'?��I͟�ϧbB]3�kS��yc��Zy��Ԣ����z�I��_��S���'�v�T��91
����]�s�"Q:�o�+q,���e��j�֧���ʍ:�2]b�M�*>�@�wDI�V�҄���'�r����f�OB����Hp��� &��Gy�iD"O�� ��x,@���+8]�ɢu቎�HO�S$X�0�Ѯ)em���D�!qk�|�	�$����M;��?a�����O�^��������/�LD��ǈ����D�*9�}⨙�cz�����9T\�UK�nL;�~BIY���>y��ϗa��MY�OǥJ$�1�a�e?�l�۟|��6ekB}�� ��i�Qw��i�FC�I�yT�����א_h� h�H�K|&9a����(x�͒�4z�$Xz�� I��m��ɨZ��!���?Q�����O��Dy>�,�O��؉q%hHpq.�Wy�(�G���n�|Ұ���'.j�&H s�y*FcS}��yr�N�q��ȟ�j�	6*<50�E�dB�M3D�(pǌ�����b����ԑ�6j1D��
�]��zA��dQ�����n� +�}B'Y�Nʈ7m�Ov���|�fa��`���6J�<��� �<i��?���S��L(%f�Qlɧ�I�>6����IBXy���n�cwQ�<y��#tlxD����7������	2�:pk�,���(O�����'���'��\>���?	��#����8�3u�����?E��'�R-/U@��󲀞� CI�Tn�}���M<qf�=T�嘏�����<Q&h�1ћ��'������'���'�pl��h��K
�p��Pc(�����_���T>#<!%%
<�J�j���%� M"@�R| ����O"�1f�	]p)3+T��-Z�"�1c��6�)��T"��?}(�0R�T�0��(�E"D���q-�=H�P3�S�R��Uӆ�=�%���'pb�`v���[��T����C�v�����?�RiҤk�f�'���'C�I��݄�������#Y�$
0�ջ��	4z����� ��g �)��̓�fM0wƘY��O���f�'��Z���Q�`��I�!��E�'B�������=1��B�i-̬�ײ���ȷ
N\�<�GH�\P�SL�J�t��I�5���"|B�bϗK��� (Q$ָ��Ka0�0�fV%mb�')RP���	ϟ$ͧ/U�<��ٟ$����,�0�BGʦ,@,���+(�O<��cX����O���p��$�#-���1.$�O��;0�'?2�O4���z���5d�H�7���y�� 6<Hes���.��ł7M�y�g^ �"qH �
�WXRXʳ����yR�-���Al�xߴ�?����i�|�\�yu�Y�V�AB̚)}c��O��d�O������OHb�ʧ	R�)� �	2\�T��L�!�� Ey-���j��b��VH��X$&�:!��#8b�d:ڧ^rp9��Q�z�2]�pN������8nnb7s�@y��ע�����	<��}ꁛ%�E4��a���k$2�ϓC_Ҙ��?Q�����?���?������9e�N�A�,��Y��d_؟��<��O���I�J�J�c2L�%J�:E.��x�0"<E���:�x,X�$W4��e����ǂ�?���?�����R��U��T�W��&��l��7�y�'�}�c
l*�6��s������ĝ�O aGz�O<� 
��h�	��EЦ!�)�`+B�'��� Mj� ���O2��<���?9�J,�� CT	u��=��l?���"��2�[��<���ԣ&AX�3�K�4*nH�6�����`U��=9&H�)9��)a�%^!�?�b���?���?�gy��'��p�J ���]�8!Y��"]C�0m�l�`[�2�"�R���yy��(���?�'VqCl{��#D);��I��@<� ���A��?���?Q(Oh�$�O��S��>���O*���	}�D9��\./�`��'�bԁ(O�i�*��8�X!͎mE���'<�!P��?)@�ǩr� ���Ą�Q. u�RJ�<�ӧ�8.��!��-_�t �0���O�<Y`
T2dw�Ҧ��n�b@ ��<����S?�j$nZ�����A�d����r�]�A���T�ߗ�yb�'���'�p�X"�'�1O�ӑm.�a�+�H��(�kԖ@<�<1�F�H�O.�܉�.��C?ܪ�#ۮ=���3��$<*R�� 񈩋� τ����J��Y��C䉿|.����(w"�{dMPk���L�;auEQ"��'/ٰ5NǄ�d�I�t6�r�4�?����䧝?���?��eɻ`�Z@�7*@��x�� J=sT|"������I����L�`s��I
V��	�	�B����2NM7�ڝA��,8v��B�n]�z���pc�'���)6�����!ј�dL:e��g�>�S��z����gx�xs7ȕ�Nk1���
9�V8x)���D�d�9%ۗ&��(��@&M���?�'+
���'�r�'��������	�f$�A�ڣ,d"�!pၵw�N�	�u����
^���.R�L���kb�F*O���A��}¦�r�b�#Bi�P�$Qsp���~bK�?��-����G�X�ғ�:v�6h�ȓ�L���
	u� e����9CP���)��<ٵh�2Z�d�BZRUsQ�<Q��M=L1ЄYqg�|O����t�<q���[����B\5uE�E�4�X�<y�Ï*$d�n�- �$���nMQ�<Qǌҗ$`�}�)_(#�V�H�N�<9�+��sh�h]���8�B��M�<�5^g���E�V�
�P�`�o�<iC,�1NH1���%@z��(�d�c�<	� ݸx�\i�ǭàu��i���a�<�f*B��a�͗x)tdF$�]�<�����od�X�Pk6izX��a�Y�<�&�J>Hꑙ����)"@`QO�}�<I��
�s��!��5���Ku�DO�<A�S�?)�J&�;v{\]#SOVL�<� �$��MB�[�X�A�Y�.-����"O 8B��6��,�ÏGp �"O��s�)��K�p�*�N�.ԕ��"O�G�5�8-���	�c�M��"O�A��2�D�[���KP!"O�tj�6e�J�A2n�.U��m��"O�a��.�(s*�
UO��Y�"O����w��� " ,�0�# "O��`^�@6N�Y�-ƕ~��Pj�"O�eb3�
���S,G�GN�|� "O����)Fj�)���R"O`e�Ƌ?�a1�$ϲo�H��S"O�;w�
�K���´鏩�b�g"O.�5�0�"3i�=7�^Mؕ"O❰ �Y����J�|�$��"O�����H+��i�Ip]���6"Ove�|�%�'�XO�*�"O��S�B�"dn�)8&�;(g 	�d"OB����q�΀�v���W�t�"O�-Z���* ���VjJ�"O��#��
�X1��J�xF��"O��S�f-Thd:�)ٯF�)Q`"OX,�i�.M����A�<��u��"OB� p�|q���o3�i3T"O@�)ciUȌ�J�H�y�9"OB��r�H��$U1l�<u"O^u$�m܊���l�{6��Z�"O6���շ�������0�4�U"O�f#и<%V�s%*.�X�"O����B�F�������dm�3"O� �ݔJ�xHG/Ҭk�0da"OfQ����K�X�[���,��DSG"OȨ:sE�8\U���΢}�T�YG"OP�g��
y�TJBmsui "O������h����TZ�l8�"O���G�*����R�E#?0HD�"O��A ��t,���Pn�w9Z�b3"O6�eh_�ߢ�{A2p���rT"O�-[��]�!�'��Z�ȴkG"O�w���l[�����O�P5��"O����)��VŔ����S�=7���'C.��K�0�D�[�H
8�0bg�.�#��!D����h��Dl�m����d��
�@"��5]�h�ᓌU�4Ta�V�by �eڧl� B�I�Dx@9��iPH9+��=%F��
ā&��z��~��\�16�x۱���E��Q#OȂ�y2��(g�`��EV�5a��Ԉ�?�����0?aTj^�`$�;��Bk�2�1l�H�����+l~�	��"�h��	�56xq�����yd�=x����M&?��[b�M���'Cܕi��O����=��	v������uR�L�e��%0�B�	,r4��R.�r
Řu�p^�b�Ab�(#�HA�g��s�\2	^�j*d�AV P�2jX�`�2D����<S�� 0�@�S:M��b<�I��:L���'�J�x�RR��)�'�L�{N��	�'PJ�zT�1z��ڧ�ʸn��I�b���@��+�hYH�E�/
A&I�`
M3U�����I2m"~P
6�d1O��E��Ը�(󉏦#!�ӱx�E�uG�:�j��#HU����z���8e��0�f�
@vq�b\kLB�I�M� #�D�8�1�	%Xb�赀0P��O0C�������H���薨]��Qؐ�E)X'!���/�r��h�[��,��>B��C� *��' � a�����`[���o��U�C�6ⶢ<�%f��Ns�aY���/!�T�G���� �uk !ܔr��\���q/^т��J�B��lk�F�5Y�����hm�uE~2
K�Q2�% w��xUz�e'X>#�!kO"�O�j����$���s����V+.?�ܯ$��rਊ�k�RYi�n�)_��H�@O��l�1k��Gf��HI&LDd�B�Ķ_3V�dF�A�7��h]x�S�$*K5��Ή�� h����=G����i�9*a|Ҭ�����R��ߪY\��`�H�3�*�H��Ar�j5�K>I��Q?�?����H���:W��h�Q�������v� �ǡ�̝2�#;�!$fNꕅ\XP��WN%��O�P�%�s�4�(u�4P�p�%�'�2q:�B����B-�b�R��dU���.�/�X������`CR���Amb� 􄕸=_|���|��e��KżK̢��R�xB�˳K��p?)G�[���!��$đ�'Ypx���#I�2�0�U�#�ZD��NM�OZdk�j�M��ly�.�F��4y1ɖ�"ؐA�-�%
h�uAa�=U��X�k3ړ�DyIa�::�P���L_5q���o�㐆1[�� "�wY^��>I$�M�W�<��7�S:FDl�Y�Fh≸IA� S6.,	묌k�`W��$��%cB����ژ�v4��C��	�Q���3���� ��עp�����|�PZĂ�H=p,�9LO���"�D�O�6]�W�K!=<F��% Y�lBJu���w�<�"Fݍd��Yp�Nn�<\��I6.W<]y�ƃ�Q�,@BX)-�44���`}F1�鉶�	�V�H�~#��蔾Ё��B=98"������P ��;�/�`%�TG�Hj�xC�-QT@����*�=��+��U%��v`_�Zޤ�<�rhO��ޥ�f��3<��ZQJ�I̓MB��Bv,_ $�&��B�M���		$G�BFb�l�إ3�)^��>)n
7D5�x!��h�y�nV�ra�qAPk�� �2 �E�ֻ��<A���7i�x1&2Ba���>L|��'�O:9�f��z��Lɒ��"��5(Q�#�OPLiT�^'GR�yʶ�]-Q�� эC.v�8h��'LO ���)��4u��C�%o��c�l�8GڼEiFO�+_�2�r�� eX04Ɓ/њ�Q��ǅL6��	�8o�=���ս+���e�44|�O��m�[�l1�wn�h|\ܹ����"��y��YrƄw�b����"C��Y�I�e�`MzC'F�\�!0���%9K�>���O��Š�N��[D�!w%&?�~��GM.:kd��A�!?��!���O������C��A���*ZB �e�)
�^�:���Qjҽ*)�j�"�,�xpD)O���" o�'3X�!�9�5ؗC��D����B�*���'J����ITL��E��0�]s��Ͻdq�	peϼ�ē;I�r�'�(C.R�+�r��O����+�|��%��K��R�;��|DxroʼK�<�4��y���*υ�M�O�z�1��V7d��a+6	��?1���d�	�iv����`��x�'����G�2#��xB6j�'l��@ǐ(9�)1栛$#�}�2$@��M��اu7&
��Š�RF����~㢁��@l8��]c��{ԣդ?����O��uU��	���k�_�)�)�(k���dĀ�
 �Q@mˋ>�RC�����a'�,���{�A� �8ET����&�d�J��� �J���i�4[,<�@쟇�V���IC�-I�'�L�0��'Nh�Pr�Z�G\�Ժv����D*c��!��x��Y�+��y�\�9��JɁ�~�O(�e)�!�bl 7$��������h=K�O���"	�&j\�p��ǃ7&$�C�F�j`Ip$�o}"a8*��Uќ'�x�����;���+f���*v�ΝFr��p��(Ģ��ϟBz��0A�hD��`r�*xPp�q���Kބ���ѻk1��@�7Z��D�O�����t��V=��'��٘u�Z�g��̨"�{XfLCI>��Pvl������{r`جj�Pฃm�"�R6zb��ai���3��(d�'�� c�hX�`�f�Jtj8��U�7n������n���C��*�Px�§\u<a�b�Z~y��2���Z�b�qF��c����`D�=L٣	�'b�d��������n�f�^̑A�Z��,9�a1?�'�����ǧ4�5���Oj &��*$
��XC�����QLwx��È���(�UD"��еM��{�J���a�9H�d��#@n����(��-���	Q
�/N��@$���4O��s/�Q��I/G�(`�:�I-C� G�	s�H8�J�0U؜�p @�"6���	�:�U�	ߖC�nE vD[-Ş��J�.�l;p�F$ ǴԄ�I�vmݛ!W{����6)�-I�\��,98"���^�	�nH��"N�v�=���Iq-BX�P�X?�,yɇ�[���x��אdw^d�E�-|����m���~Kr�U������踧��D/�4�λ8�`�ц��:{�����"��A���xO`�CcL�`�b�`�0G��e
 d�l�N26n:[�2����E��8$�p���0{�J��s& Lf.�BA!O��qR�V�s� `0w�
H�8I��흎�����X�0}� �'�芕���9���	�/Q)R�"��J}�ͩ�	�H�}	�����	2'����d��P�'�y4 s�'!�c]"����N�)�z�K%�9U�Y��S�? �q�C��V��z�m�8ub,a$�9<��!� �G]��S�'1j��'E��s�BܻK����/�cw.�Z
�'w�9��WRz~(Z��*P2��J��<a%熠q�� �)S0+4��$��)��y�'J�\\$SeFL� gaz=O��r�&@B?�Ң�Q�����ڼq��i�@�`�<db�9 ���j3�FO2��wB�^�'/$�Q�b�{�Oj��k%,XRf����56+�'����r����������Bl�e	.-<I�'��Ÿ�bRm�g��*r|�Qہ+Y'�%���Ѐt�XC�	;:�%�� ��tQ��;a˅|ϨlC�O[0H�i�%���p>!����	>�pF ��S2�ʄ��u��A8I3�D&�8�D��Ov6-V$���]/l�	����T�ۇ�[�>0!���	���U�'���y �Z)j�J>����{!����&o��M�'9�N�Ӑmʓe�T0*���-�G/��)��B2W�Bi�.��E�P�"�Bޜ�Mf���ы��M���L<Q��F����%�<?Ħ�*ǉ�w8����N�4�1O���#W!bt]�vh�9s��,	r"O�
�&�R�@h��fA�O�n�7�x��̀>�$c�b?ي��$��q�4⇡J	�#!?D�`�Q���.�XM�HHŪG�;D��(�)�[L�Gg\).�����9D�h
�/HRP9sF`;_ ���ek;D��8 +�\��LڄF۶*�����9D��K@o�	2Lhj##M9y�hⷀ8D�dR7���k�5��a���D]it8D��#�J��r���?#Y�<�k7D��R+]!BY���,�0���F#8D���曰J&����P/6�ܠ�(D����_�GhL}�0�P��$YPD&D�a�aV!��i��B 4If�S�F"D�T�)�?s!��zP�˦;LJ���l D��Cƚ.�$1��Huo:��f�?D��Z���<  Y	t+Śl5(�(D��Ⴣ"}X��!g$ZI@�(D�����S�f��1��K�>]#�g&D���e��L���;�k&�d�!K$D����M�$��� ��H_d	��5D��(����\�2����՘|z�j8D���	z��4�fФwt�1��5D��rQ�1@g:m�@�1�&hY�m2D�x;a�4h72��I�J�L��e%D�T�GڿM��lHc,�%FQn(���#D�ifK�7 Y�Q �� M.8��o-D��肬�+j��$(� :RA,�jfa>D�0��H��Rő�ė�,3*�HW�>D�Q%H/k��`�F�I�e��0As�7D���b���
��i�qA4aA� ˥k+D��b�ۺ�(!j�MZr@��Ua)D��P�`ӯ�u:2�)����C&D����!t�v]8������� �%D���
��4DP�F8q�$��H�<yD���*��0"\*/p����Y�<��@ܲf�6�
�������@�<I�ݡ�1"w�N!6�ΐQ�I�|�<�%�n�v�r#�H44H!"Mn�<F&�&.n]c��?n��)�.�t�<��F1
oHg)�=Z}}y�/�|�<���̠1y��%��m����z�<��@�\�d.�5_��D{�\�<�DfP9Y�v�%+��m�����m�<%��06��MiS�U"��P@R �`�<�j�$N�hr�� k q2&HC�<aX�`����@Y��IJ��@�<)ׅQh���cM�h�jM�D�{�<� �D�p�"5�sh�|����"Ot�����h�t�i�&�?b�x�"O�m�ĉX2{�6	��B�J,8�K�"O�ek���Ms�I����/zr,+�"O@���ÍS��l�&�Ėy�X�@v"O��+aa�i��DKD�_"�N�@"O~y�-��0����B�l���"O�hs�d/p�������4��Y��"Ozh3q�حk�b�Ro]+ٲ��@"OH���m c��Ġ�-O�i���#�"O*�:��וt�TIyو%���Y�+D��`,�X���gW�w0��ch3D��@f�Y+hK�᣶ԓS��#+2D��7��o�V)�GN�"v96P-4D� ���un �!I�!6q p2�?D�ԲsB�n���� �֤��	J�d!D��"E� #��C�!J
TV���:D��!˛�lPH9����j��h9D��xa�N�2ɘ�I#E w6�%Ag�1D�TiƎ��U9�Lh�I��#U����<D�l��"^>V�����@1\+�Q��.D� �I^�g���ue���bw&8D�P���)R1���g' �\��\!�)2D��r�L��Iޘ�pu)�`��B�4D�Lâ��5C[���p�Y����b2D�D#5).��`raE�5<��(QJ+D��peǄ��!*����1��*D�4��`��S�!ܔ<���R�-D�@�K�sU"�B��
Q�+\	zS!��i���)H?��!���τ-O!�K38y$��7�к-��`��wF!��ځ}�0����,(j����"eL!��sZ��j��jRܣa`ʹ}Q!�:>�� s����O��y��	lF!�Dߔ77Tѓ0ˈ����@.��C!��[�N�s��^.Mh��vk�3!�Ē>�BA��H%S�Z�H`�.\!�$ؙ#T�4#���d\��i>I!�O�D�^i:�jU�]�^��7��!�8)�FH�a%ЕN����|�!�$F�f�RL�g��<y���sJپ�!�d�"\�l*���d����/��\�!�$5y���P�Ҷp$��u�
S�!��0@0�h!��.�s�̓�Kt!�dԉ(�T@�";��R�l)-d!�DJS"��K׀Z	Fю)Qrɗ�~L!��%%1|��E�`��Io�>H!���TL�Cv� ����ƭ�TX!��;;�.P1,��NL�$��fC!���_~�P
�"�3~6�(��
�?�!�żY��cg��$mQr]�t��US!�d�)xR�3��1ڈQ3� �d*!��Y��X�ĭK�,*�e�q��,!�d �lV�}�ь��Zd��w�x!�$�1N� ����G8%�ݐ�+T�!�$ڶkCdE�U�ç{�ݑeзxg!�d٪.rH困{�l�r�D)
Z!��K�`���jz�t�q��!򤃕b����"h�L[�YcH�;A�!�D@��,��Ƿ%���q��:�!�dǽC���5*˨`ɔ��g�9W�!��1��p�䧄�
�h*d&�b�!�$@��JL�@NA)D�Q�d�r!��[��q��;Jޮ��r#�;[!�� e9�ɪ�X�q`��Z �Y�"O�t�(���� �ɓul�i�"Ob"��'s���і��	l��ұ"O�0Z��W�T�H�E�\NSq�"O^e��l]
�q@Z.>P���"O�<��j��^��xt�ǶzPPE���:�S�@�l�sb̊KT�ʁ��q�B�I<r�4D������@B�-�8�B�Ɂb8N����Y;�:���
]��C�I�_*N0Hd�_��� �|�����>)!̓C��c�S2,�ʼ��%�|��p=1`�S�j94�J�A
 ,�����~�<q���rrl��Fj�dúa �GU�<y��βa�Ԥ`�-�D��Q� �S�<����s�4ŨS+�L�@�0�R�<��)�M
�2p�ʤ`�л�d�<id�˥�h̪�M��GR�����Jz�<�cța�bZj�X�'�4��C�I�#�	�f�θA*܄ ��ܣQ��C�	�s����i_�SŬ�*�.YPO�C�	�3Ȥ�X�CW�9Ή�c،D{�C�	5Rr.���ݾkLb�+�(ęBu�C��	a'�����$4(U��C�6��C�I�W����S��zL��[3c@�+1�C�ɇ;;L��2E�[>� �G�ߞ&�pC�I�w��<��N9�|pi�['j݀B�	#>xz��c��u�B�p��C�=pB�I��}��n�6�2������NB�ɖ@�&Ip1��|�p�""�[	Z�vC�I2N��ŸVG	��>@�4�]0n�DC�I�9�ܱz� ���@A�cA1d>vB�	# �Q�Dj["(:�4��Hd:B�I�`v�A�EK�J�v��w���<'B�'�$`��ǜ�7�`Rfٮ3�<C�ɰq�,ը���^�H���?�>�IN��@�+���^ ��茬v�,�2�<D�D�0�V�h]S�
&�PX/D���b�_�8��-�T) �40��I2D��s�Ѕd6�M��n:S����/D�h a��F�B���O�,���To,D��X��$GEy�C�'q��#R�'D���I�[q��c� �*b͖ya��9D�0zW��&����I�&�8��f)6D�����@#8S�Q nI�~��pj�#0D�8��!
�x��V^���"�C���y"�ѯ�h$a���$; D��G;�O�=�OT�%ғ���{��d����[L^q*�'5��VMN	;�J'�ϊU�D� �'oz�pP��0�X�Q(�-N����'#d���)�!��X�����>����'�^L�$h��uW��j�9$(�E����'xȉ�6��+,��ВL�2�$E��'m����Ǫn.��bH�}.0��'�.�v�˱�d�nА;�.D "O�ѱ5�U Y+��葯Dr�Q�1"On�+��NkfYZ�.F�G=U"O&e[�(�7%0	{1+^b�! "O� *�iL�Kw���"�a��e�R�'��IG�x+�c(f��Yٖ#^86�C� ����"EƆ�#p!���C�ɾ@T��iF _�p�!���M=�C�I#�̸��m��O�h;�/�Bjc���'WD�~�" @	����)�	Hް�*娔g�<��FNW(1;6�ۆy�|��$�<� ��P��/y[PT p � h(�J�"O�l#���'����1Y��q�"O�窆�}DP4�.[8(W���"O�4Iю\7Ba�Ya339��}�"Ot�6f]�@�H��AU�|:l�"Oޥ"f�W��Zl�BK�:^��#�"O(��G�/V���놹�}yP"O���4��@tÅ�_	�����"O��sQ<*�R�Y1��B.�%"OH����IRf2A�>K�:�z�"O�����K?��	��aСJ�"$��"O�A@�w�P`a���b�"O���H-SJ��EJ�\ؒ"O���J�}t�(XQh�-/0��"O�U��	�f%�0ABB�<?R}*��x�E[���O��	C�K�9 � ���K�H%X�'�p��V��Jw x�� �[B �R�"+�eX��@���'}�
	WoA	O:h�ע<D��i�W�NI��B&�_P�`�e�Xh<�UD�>���Z�e΂R�n��R�<�GCԔ�T)u!��Y҄���FK�<��l��f�F���)%�5��BFL�<)�T DgT�d�@�3��}�&�K�<i`lз�@D�c�J�j=��@�@�<Q�ܨSf<PBn��!֬��B�|�<���#4�(�)�.Lz����@JNA�<��G'k����b�#VQӌQe�<��-�ͅ�J������*05pa��c�$R�"ġg���a�T�[��ȓn��I!�/�X"� �`�0����ȓAFбѓ� �N2�b.A֊	�ȓx�V�z�&��C�a�w�ͦ���ȓ2�3��1d6�'�#��ȓ-�.5�-�31ND�@��!�i��	�����MC1cM��Б ��j�1�ȓ#!��3��R�\�+����ޥ���O�Y��Rp AxE�,D���u���^uTI�7E�*�Ҭ���5D����G�8VXQ�'�P +~~�P�%4D����0~o��H�,k2|H�F�3D���t(Y7�l̩Ċ͹�X��Aj6D��6d�'|0|��a���4���5D�졥�^��x�	�LԢ	�*䘓�2D��x�B;Una"0��
����h>D�dX�@��M��-W:k|�M���b�<�0��?���Y�0�r��D�_�O2�B�I��R�zP�V�;Li1cb ��B�aX6�9���.�x��W@HB�ɺ0�@�M+3�����	;B�	,�\����)Oإ�$PD��C�I3�����"�?]�D����ZC�I�hѻ��Ӗyn�ѣ���CA�C�I�f��J��ۋ ���cC��?H��C�ɼWo�hqa!e����Fی��C剌	��p�.؉d����f�
d]!�D��~�D\SGǹ~֬�ehN*hP!�$��0^�� ��hł�
���0P!�1� �`P��W�2��mH�^!�dZ�%��9�f�ܡx�h��i٘�!�	0���-�+�����"K�j�!�D�-"\��AD�t瀠y�$���!�&c�V8�gm܄O�&�xEcٕI�!���_��Y�E_�G�6�CW9I�!�$��t*��4�ӕV��9`��Y/�!�� :��GʜC��X ��<o����"O�4��e��X�x�H�&Rb����"OFX�#Z�"2��U�-3|��"O��r�ϕWl�1��Ȉ�7"O�| ��N�N@��L
X��%"O�	������U��5/���Q�"Oz&jT��ڱ˴�[�M3�:A"O���l�l)pqA�.� �
w"O��A�EɃ	�|q��ޚ^�rl��"O�P1o҄*�2��#�;�LmZ�"OЕh�/S2!�4Bǂ�Qy�,��"OM�*L�1��a�t��Wg|��T"O�̈G��M��c��hU@��"O�P�C`�9����rk�	Bۼ�;�"O�5#G��G�^r��ڮt��'�v�c5��m[)*!�N�f�pP�'0�M0�)\�/Th����,2�z���',z�2DƁ:2-�<:�W!&�ZI��'���I�[78�~��B��%
���'��t��o�4?^�8�)�#�	��'"��Q��ah�jQ'ͭ�bpZ�'���2�W&��<�0'�!7Dc�'w�`�@��SE`9+"��5�A(�'��Q���:k������X:+���'R��p��W	�Ȱ��ʢyrp�K
�'��d��нm[P<�E�ȵi�0{�'�b� &d՞<<X���Kb� ȹ
�'�nm#΋�%xP(c�#��]Z���'��b	�8C�*�KٌT$��;�'ۈ�8�(P���dM׭6�l1��'��k#�]5{#*�@͈�/b����'���*%����ZЃF托�T��	�'�.X*C��r3�]S-�/�a	�'%4U"��')��[֌�2��j�'F �����<��i��U�~t��
�'��Mdhw} �!�Lmq~$	
�'ena�q��,�T���T�nW,�	�'��H��
�75�^d��T.j����']�\�PGA4/U �O�+�)�'�\������~Y(�ڭ%[\�!�'~aP�f�?�RQ:$@���lu��'=|�Y�!< <�C-C�9����'�p$�nK1F��3@Ɖ.�N��'�⼡�I�d���"IS��
�'�vUc'��/DHh<0���[��z�'Vi��@����喂|ԡ��'\�)�#X0�R!C�w���'k��{���3d��T�bE4���'�؀9S��~�Ȱ#��_٠�(�'a&�c�v�`�B<Yx����'���
1l'M� ��Z�V��x�'�����ߏ{�@3�	�k�d��'��;�أs�H�䌒��P����>P�� �d���H�e%*�y2��,�Lʓ���{$�L��!�y�����```蚔u��@k���ycT�	�����f՛��=�e���yBB��J\�U���"r�T�رF��y����|5`�F��n�l�a��7�y���+L̰ܩ���k�ʥ��Y�ya�8-"|�aBHu�⡠'��y��ϓ�P�QDG�; Pu�vI��yBm@$b��W���xQr]�6  ��y�X�/ծ��#�B s���+���y
� v|H�@�!r����Μ%x�TɰP"Oxy#���;��I'E�5���X�"O� 9`��%cc�H����Zq"OL܃bװll��uF%0���1"O.����Ԓ6Z �I�Ĳ���"O�)RK&SMP�{��T2�r`�u"O�`{1N؞#y�D���sx�e3"O�ȠW���I�֠��g\�i�"O��3f,;IjA��.�"5M�ܫ�"O�0��E��X��c�8]7�
"OJ�A���_�2h��(�F1����"O8�ËФ�4ݫ�h�6���1"Ot5��ޕ\��HPH�1����"O*�rA��z7:,������-@�"OHI���˲u:����m�\�"O���c�-0��Dr���?�ȹ��*O�ua��� ��VaͪgN���
�'��K3M�~�|���	�%U�L={
�'2ęf�J.���#B�X�!��'Ҩ�Q��8j���#��.I���'��m�� A-p�e`�έ@C,��'$x �Y4K]��B`Ĉ@m����'R6�AQ`ϊGv0�0�Ií<�vLA�'���vj�C�:�Q��� �%��'���сD( �ޔQ�.��"���'|i1�f��=7�ec�^�}���'/d�j�ĸG�Mxt�Ov�(��'��dD
�8)�t��*��=�����'�j= 1gC�W�3�/[�Z�'���5��Qb:�9����q$!�'�V�qAд!:��;o���
�'[<	y�Hջ"��� BgZ`�!	�'��ݺLM�d�@AwM���ls�'���0	ҧ*�lPfʔ�m��
�'��\��>N��0�� �)����'m	���__0`�ǃ�-����'�~��#�2e�V���( ��'��0��"X3}d�4�$�l��'_xt(�f�0�8���D���'�$���3qQD�iшyb����'��zv�ǁY����!G_'\�^���'���Sf���B�	��I.l�9�'%�����D0H�&�8aA���9�	�'�(:v�G�H��5�4KΠR	�'��� ả=[B������ygZ��	�'p�`�Bϓq��!鳈����8i	�'��ȠѦ�
�� Vg�>�� 
�'�2%R�$F*� �� �T��	�'爤95�B�l�
e[E)U1����'ڤ�t�E� /�aK��4;Nz(�'>����l��C4s�H�=8a( X�'E�D�7
݈$��mz#K�)�x�
�'^p&��}����d!	�AP	�'�"�8r/�<�����
� ��e��'O`���b�-VvAB�-
�^f\��'arȋq�G����Q@�����'�H	�cO8QXZ<Q�߇#s�Y��'�ā����hH{�.��܈
�'������Z�`��p	���n\�� �'��D�Q��2���V%ƣc!Z�y�'�k�&��)�AKU�	.�T��'4T��p`\=9NiCI
�'g*���'��Iw�]�GV813'��.=h,��'����tȞ	2]~Q�특��!Y��� $��0��)
zTȳ�͝;|���1"Ov��'�2�NC�M�|%VyI�"OT�⠨��idX �GA�ػ�"O���T 9���)AN1X@�"O���"���LĈr���E$�Y"Oxū� (g}6����M�2"O���҆L�~����ϛ2��E"O�0�&��(��6M�V�08P�"OZHQ�ect�Qv�ƧW����"O�(s�@N.J�<�����N���(�"O�)ȲO5�T���ÃO���'"O�Qc��6UCɂ��E�5�����"O�����W'�	�L_�~r��7*O�1XEF���P�5�F�}V�X
�'���S���7Gj�+׀ä-y	�'&��U���E��1e��z�ZA��'.X�ѷmȦ�ޅ8�瑭Fa�{	�'?j����Z6t�O�>(�Y:	�'lE�`�R6&�<���90D���'C0h��J��Z0���{�N�9�'U0�+����|�0�k�!
���
�'���тh�%_�%z��U�m~�M�	�'�q˔���UPtq�잏b4�y	�'4�U��+Y+�&�0��B7P�vl�'� ���/�'I��A�"V�,j���'�4�d�HL��T�^�P�'�n��5Jۉ�����DU�T5*�'�f=y��0|�m���1�6���'�X��F��Ӥ��4��,��'�4�6ʁ,!� X��B���pY��'5���'"��G'/^v�A�'}~�x` ��TYN-�d�TS2���'s�<��HQ 	sy����L��	�����qy�,���_�+�f4s��U��y����'D���+"��q)7*_��y�E +d��"t��$.Rx��V�N��y��(��)��Ӷ&HΉ����yB���x��9d�^"$�|�����y�ˍvʴ܂v@��"B���_�yB�CM"�d"j��q	��ɝ�y2��$�
�)���*���y��E)Nݒ��E�
}�ȀO��y�ڶȼA����zf]�P��6�yҎ�4f��8X�/D,E��G����y�Q�4���$�8X`d�0�y@}��@�u�R|�2�M+0�Y��F���C ��,6���@��R �5�ȓ��9ZC�ɣ�%/�U[ m@�"Oؠ�U��m�$!�nC�kwj\�F"O, �������#�`�U��"OƜ��$##�L1IH�`J&�a"O��Y�d�1>�lQ#�Y��α��"O8��Ƙ�!tNu��+�~�f"O��d���;.t��+i	n�<�y��K���i�(*�A&bZ�yB��;%"ܹ�n2�V��J���y��&����$��FqUb˴�yr����X�k��>�j�d��+�y��M��:�*�`��hۄ]P��.�y�-��
_�Hshٮe	.m�&�B�y�H�1ȹ(�홣���*�+�y�h̕pT����};�X
� �5�y�F
{� 	��d̜>PV�;D�X2�yҋ�5H�<�#^N�,"��F��y
� ���/�f���`G"g�ۡ"O��T�f8`h�A	�i:�T"1"O��z�B�57���������2`"O�A�@�4��2���m�t	;&"OH���݌^�~x%�"
q�A��"Ojx�#� ���S�K�*&mE"O����L�w��qj��pK���y2�G�8���jнI�\��� ���#�S�O�А#���u��� cč�+�i!�' ��ⴉ�,	.N��2C�)�5�
�'x@m�S�:S�7��7$e"�"O"�x�cڿ%I�)��W8J-�l�"O�m���*���"$	ӹuG�ԑ"O�UڔE�;87ZA����^�]��"O���� ɀyb�A�V��tO�f!�d��`D��φ2d��i��.�3.!�dͰ;u A���<$߬��q蓩q)!򤙔��!pK8x�,Tq2�ɟ|!������@5my��1C���4y!򤇤�"a�%�V�~w����h! "O2�ū��nV�EȱeيM��I�"O$8��>t��p%R1]���E"O^��`R�2#дS�Fűs�<��A"Or���`%:���$�1,j��`Q"O�U�e� IRt�bѾ2J`�"1"O��RӇ
E��HT��u�&Y��"O�-6*�7,��aB�d�6$r�"O&�#��ěC��i�A�֠2�O�⛲?
���&�)j ��B5��<a���'E�(��ǀ�+�)h��
?�t��M-D��bgfB'<u�y*@�	�U[��B��)D��9�F�,P~A�fM��D���-D������j?.TZBO�c����0D��qA�3,�9�j�a7�Ak�.D��:��A� ��	ǇM22-����'D��Y�M�y��M���G���GI0D�dh�&Cu�������s�pA�N D��ʦ�+�&��eJ=g��ڠ�1D�4`�̜i��K��Z.U����g�+D�؛'�R#'4H���FY�O� �F.D�P�#ă�2�E©�)B���4�*D��To��%�]!�H��A�jh@.D������ivN��ԵVv|E��E1D�����׷o�8;'W�0;B�Fl,D���N���Qg�"��<*��:GI!�3�� 	��^1z��d���э<!�M�FZ" A�gK�����bu�!�� �O�8l[���O���į�b�!��@�<QFDK�L!���HWe!��A�Mxv삵M�xtB�pE"O�B����-4`���1"!���"O�}+��VHm3��ݻ[� �9`"O<��D��6c|�PD#F�'+4���"O�}�p,X�l�E��Q�&lh[�"O�H�UA��VO�ٱ#KŽc�Z,��"O�e�"�DK䫂D�8��ĘW"O���eF��V�!v���p�4"O���fŝcZ6y"��J@`��"Ot��)�	U�"�0)@�U1��ˣ"O��r�i������蒙P��X�e"O��b KH*���QW���s�E""O����eI o/�H�3��)[�a�"O��.�']��u�E��vX�B"OZ����_�j�Y��[�qr�%��'3����O�? ����'ȝK� `����&xhm@�"O�تa���T�*�@�ےiv���"O���ӺyP��q��)lb�h�d"Odً�C��1Ԉ9ԧ��]���"O�1�J_�-�g�"�d8s"O
�x7%���xt�^%1��L g"OT@CWg�N���P��(h�`ⷓ|r�'"^�J�p��;�[�[���!
�'��U�lZK$y�T�PW���p	�'~���/^� �0x�!��!&P`9	�'�@e��=N^�1� B�<���'d*�d�6nN����(5���'8j�*�k
1����M)D����'��E�Ơ^-��i�%�=��H���'x�i{� �_цt�� ��>��'G�q�bԌ�pd��ˆ7H�M�'�>4����;�ސ+�O��0��	�'��{���U��B�ލtc&�	�'�BaVj�*gQ�]� �*s2q��'y��Pa�95)�xI���q�Z�Y�'2Ҹ+Q˝�!|,jࢀo�v%��'��A;D�#O[��Ⴃ[ v����'(L�A�͙,��,��%f�nYH	�'����1��C�0�&l�RT���'���	��vY�0�R��"2U�!�
�'̾2GM/h�ٛ���\�֔�	�'(�@��5X���eۈxp�x	�'ʲ�`���'�lY����Yc,HC�'�����3�� f&��G��-y�'�l�y��ҟA4Z5-ľ:�8�	�'�~$04��WH��D�#�e��'_XuZ4�o��BE#{��'�lX��� r�\]s@�(L�^t��'�:�0��̏f������| �  ���y��
�VA���
�xy&	7���y�"&j���q�؋r����Ʉ�y�/ Zi	���VvCY��yrQ 8�Aa�L�.��%h�y��K>-��!#V,
��z:�O���yBGZE�xT��̵���Bݖ�y�l@�3����S�b�F��ĵ�y�戻-d� �3I�u�ٹDK�+�y��B/��A	���v�f� d	���y��� o��<зjU2sX`���˦�y�@ǚ9��Q���;]Δ�5�B/�y���l��9�u�>7ʶ������y�d�Q��u���>*��]�HϢ�y�ˣ'貹�FE�
(�|�+�M�y�*�).��̋��,T%�� 5O��y��Q�"� �{f��E�z���ۛ�yR.�!7F�i�B
7|$�S����yrɇA�4!��ǵ+���B$��y��[iĝ���J��c�l�4�y⢞9}�J��4�ٮY��1uC��y��ٿP�>��%��A��t�T�N+��'�ў�O� 쑗�$A#���#��=�%��'!���O�j�6,J�>6� ���'+��[eC��YYPB�;d
 }��'��14��x0Ido�E�Xs�'E�مhW�v��]��U�s��1��'t�tK�
̘+��Hbǈgk.��	�'�j�iw�K���
OB�e���'́�o��*9B��d���_֪|��'Oj�i���g(���7nC,`�N����� L��҆
��Ƞ(ڢ2�6]Z"O�(T��
���v�*~�hA"O�����=%�A�P�D��a"O�];%�`�l���^�x��y��"O �b7��$�aJsK���5��It���4	I9� ��$4����g,D��i�'�.�8�*՝I�Nu�#�)D��(�/И����U�+K���(D�0 q*Y,�|��d U�zQ$��@*D�x�eb�` �|�Я�LT��G&D��P�Q�4��dO'��e!`M&D�Hg�W�="͑��޷>5����%��:�	g�'id�#h�7`	ZŎI1C��M��'8D�z&Cy�:���):����'`�Bf�K+x>)3�B�W��`��'���9�E�'G&M��)
/;�^�)�'=�����(��Dj�@P	4���'�8#tI��?��h%O>2j`;�'�2�	��&��h��H$/RZ���Z�x�'iў�O�>� �T�+�����63�5��'`�
� &>���%H�
�'�*��e�Z�<�B��g�hi���	�'��)�#)�)1�fM�l��g�-R	�'�j=;�`�	�J���M;
u�|A�'���ar61tZ�S�"�0�����'@b10S#��%������.�F���'�d� ��L.��|z� �)
bt��'7���kD!�*b4jJ�F ��' �eY'n�$��D���*4/���'��C��f8qY�0��
�'z�U��	��1mRdCC��>)-�!S
�'J��("M@E��f�52�e�'�4P��*l����/<���	�'�@,k E�M4m�i�w��[�'��p�@f��Nh��ゎ�&h�����'I���C���a��h����R�+�')H��Lˏ[[�������Z8�'�,�0s��R_x�Cq�Ȯ42ܭ�'�P��Qkߤ2s0*�)M�%j|���'D�)��N�!1��!��%Ϣ�s���yR/R48n��IRiͿUڴ1h�S�y���(���gҴO>�q)��U��y��-�6���M:O�I�m��y�A����,c��
FsD�X�◗�y���D��1V曹AZۢ���yR�ǉ�6�s�E". ,j�-�:�y�,ݔb6
�l�����'h�م� '�h�h��Q8�r��	�'w����"��d�����X8/�J]�	�'��]{�斓H����R#��uS�q�'ݚI��G� ,� U#�G�p:�K	�'j��  \�V��H��P�~�X�'�d8�wn�4���K�M��%0�'A�����.5\�� J�zT�
�'��F�0�r���F��o��`;�'�vL�%n̈VB�:�y�����'�f��3Nӹ#��ળ/�:?@�
�'��,c�M�e1 Rm�e��i�'(���DO�5��y�B��d�Tp�'��;Q`D�15:1i�+Z�F�̰��'�4�ӄ�]�k0�*Q �A�he(	��?��OJE
0��K�0��� �f�
Q�f"O$�PbhSp�����:�"O��P���hEhuj���"e��X!1"O� J)� R4eM�s��B�Փ�"O�	1��O�t�2�O#A��;�"Or�S`Q�A�xD�f�G�0�Lc"O
�͍5VBt[�)_�%��d"O�sNO�9" ����� �d[�"O�T"�ǌ&:�� �1�8�8�"O`�įC/V?e�C`G']F�9�"O�LA4_�l����F�߳Wހ�v"O�C�Ȇ�l��!�[2T͢1�F"Op1*"�Ł+/�<��S;J����"O$9E C5~�SL�8v^�g�|B�'g�4L���(�'���ekX�5�!��]���JP�M�)�ђK�h�!��."��E��9���{Q)E��!����E�WE>j{r9:s��0Z�!��'9���`D	� ��w�Y<n�!�$\\��*�˂�\�x�#��k�!��Ǖ}G ��a�U�1Sv� ���	�"O���*ޞs�h���c��I�� �"O�d[V�)g��{uB�+�vk'"O�� h��(��h�.Y�7�T�2"O�f�ŕo�d�c5.�R�^ 1a"O1DmKW�ũ0HTP��\��"O@`@�kƀOʢh���2Yu2LH�"Ot ���сM�H� F&�3Ei�'�IO>IIb�*Z3R-�"�! �p=H��>D��sC`ܗ{�V��t��b`}1�;D����)s����/��.�D��B:D���W��3����aX"!'ư���6D�� �A(V<dh� ".6��˓�/D�4I��@=(ψ�@�/��  D�D1q]!ɪ5{3a�
����E<�ֈ���[ET)�� ����g䕰�"O���7�ǿC;hPD�"b"O�ءGԲfL�誔E�'Q��"O��VR��`Mc��ˑ"I��i�"O��	E�b>Rl+TBˮk4�P;"O\و&�V�Hˮ����V�>Px�"O�PHGAD,m�b�� ߉O�fu2"O֔A�6�~t���Q��3"O��a-!m(�H@�@�9:��URe"Oґг(�W���r�͌s�A�p"Oظp�׺SȒK��V�rz�Y""O*��4Έ� r�y��H3ye&01"O)����2r���tŊ[kX�q�"O��i[�_�N�APDA�Gg�aHe"O��@���d��`K R�XtL��"Ol�@���9E`'`W=88��"O�M�֊_�*[���A�''�H��"O6��f�I�+��
/�-D+"0"O�`*�I�q��)�୉&<�t�"O�]��,Y���&2�D4Y�O�)�!��wT���Ґ%�py#W��Oh�=E�T9O|P�׀�N�4c�� %E2�s�"O�-
$$D=\�����̆JCxB�"O0���E����3 Ν#�P�"OVl�E��I}���E.( �\"Ou�Rą�]����L��S�>xc�"O��0���fNusUL�*T��`�"OF�2�NԂm�H����ՎP��	��IW>�����??�H�f��Jgm�3h&D�D��
�Z�$�0b�;��B�M'D�di���0k�����V7���aw�8D��hB)P�-�mה=S�\j`�7D��  �y��V)_�$�h���"�8��4"O� FV�@�4�ƋŔty�@X�"O�9����9T$@�h��çPHXY��'e�O��}��]D8��ue]$z�$ ��:d�ȓ-g"i���>U��"f 4jlx)��QV�5�'ΗRax��ѭ^m�܄ȓtO�$��EP0@�άM�`�ȓU���J�6��!��)��r����ȓ-�I �% *ɤ�JQ�!:��d���5P�'պu���!$^��ȓr���T�H�^Y*�!�M�T*���#A��x��''0ȑ�+U�s����"�ЃcO{y&�t�I�\�ȓ<J��(*�
B�䌉���0�I�ȓX��RP��>|C�,BkU6>�$���x%,�y�Օj,@�FHM65��ȓ;Ȧ�bBCK� �t
6��2Av�y�����u�O�^��Q
�.O��ȓ=����G��$j�� ��#q!��^F��c2�Y�O���{w���m��8�ȓ`���i�8�h�;"@��g� ��M��ёNб~��7Nv�8���(E�U��/E1O(X�lG8�ȓG��TK��BP7� 3 �=2���?���~23�5bހܑrIT�_(�IH�MO�<�s��m���h@%��PQc�M�<���P�J}�/G�-�����TU�<��iM�Gt���pd�qz:4xϕG�<)�½oPA;�
=iИ  RF�<��fR	�V���W;��c�PC�<�֤�/�ܳ£�|�){7�Aw��Byr�OTpx��J2�S�f<.4��'t���4���g �a��m�W�����'�\Q%���cĔ-�T�##��-��'�|4c�OG �ttϔ-��!�'�v4['�ۀL��2p�]�s"�K�'�N�� hV>G���*GB�1R�D�+�'�:UTeD�,(`M��*���HJ>���?!	çn�����jɥVz���h\")0���ȓ�j���OR} RH��A�5U�ل�{)�9���n5 �H�S(P|D{��O��Cn�S_��q��]�D�5��'��T9Tn�86�lE��(8�^��'<��EO�*]Z2|��'Z�Y
�'�%2���5�FL3M4��
�'{>哰�G,;r�)�ꍹ9��@�'=�+ѧ�y TA�I�Sܴ��'��i�M�	n�Xb h��r�"�)�d���F{X] D�~�|�[�×�y�o[�6hh�/x�$�f���y҂��kN�A�p�(k���� )�y��M���Z�c�/j$ܜ3 I8�y��S4"V�)Xt����00�yb� �m( ���d
�o{�lQ'È��y�e�0�V�F�Q<�l�Ƈ���y�A�9�tt��N��b�eCA����y��F�iY -��I�$&3�`���y�;Qq�u�C@^-�vA��h�(�y�΍�!����
�(ujh�'���y�
��>��\����2"���nF
�y�JH&Lδ!�-[�0�l�q��6�y���B���HCc�V�t��4���y�͍>�\��'�~��!dmݣ�y�5�������}b^8j0O�5�y
� �up�c�e얹��-[�?�X˔"O��C��V�t�㦆�]��Q��"O�����>Y�T�(ہ+�z�
""O��j��K�&�T��G��`"OD�u&����&C�*W�F-:�"OFH�0g1,U2��,���Ӡ"O�C������l!`ʇ��:��"O��( ���n�����1��i�"O&��"IA�ı���-[��|y*O�P�$��H��D���/@pQ��'h����])D5lh�����.V6݋�'���BhC<l��x'tJ(�
�'`����ًf��b�.�>d����
�'�yr!��j��L����n�ԁ	�'�Bt��ML���\�@5���"O�)+D���y�d�т+�x�d"O%*�N!9��jw���d�&�P"O��c�͒�MRW��m����"O�B`��#�&P��
���a"O(�j�gׁ:%�8�҄Ťx�(�pr"O0���'�yy��RbdI<|�QP@"O��"k:�BԂDd�Vh�AI�"O���v�I<o�����E1�)iq"O6���̅CT�����]#�[�"O�	#dn�W�4*� �9(��YA"Or��ō�^�4��@G= 8���'2�I.)<N(�!h޶|[��Ed�+�B�ɿT�u��R�H���c�L���C䉧LnI�	[5�M�t#�v/|B�I�|Y�ϓMPha�w��,�\�З'p�'��#;(��V� #]�(�����%{JB�I�+�҈!�Q�y���P�n`�:B�	�b�u���кJ��@�+5qNB�I:L	����$	�k�p��fӃ%�zC䉜)W&�9�K�N>Ku����>C�	��`��d.o��=3c��UqC�I7)�r�pR۬`@�M������=�
ç#��|���D)D�#!gC�q����o�"����� 7��-CƬ�8XJ1��\��Q�qbZT�ԯ^4q����I_�'trq��!�:y��]�-�d^8`�'R�tF�^�	�H�o�"c�f)#�'��cP�Ooy�IEó%�����'aݣ�n\8La��d�C�1��Ъ�'����nK�X\����(#7^r�z����$,�O�!��APh~����eV��:""O|�DV���-�u�ʷqZ���u�'����b�B{uf�p���
9�I�! :D�� e.$�� 8�-��aW�-Hc-<D����ʭnK��1�Ɖ2閱r�l6D�hI`��7}�j<d��$\�P��1�>D�dy��^�\�ăA& {�ꬂ�<D�|j4J�VNL�dѬ''����8D�8+d�U�J�� �D`^���F6�*�Ov�{r!��WT!�C�H��帄�'C�'�az�(�. �=Ѣi����g
��y�ϝ�cL`Dc�!�! I�<��B،�y�Ɨ;_���B�W�f����%���y�k؇#������bd8 ;E����x�¬A6J$B�@W$?��d
a'du!��]Vޤ�C��S�6�h�?a?�r1O�����@,�����k�Y�$A"O�y35+Q*s"p�K])K^(�3"Ov3�ж8=��ID�=�Y�0"O� -ӗ�k�
ٳ�T�H'*AH�'ў"~�@e��l��y����a�5�ը��>��OD��0�d��U!�3�Լ�%�'R1O��h�K��aE��rt*� ~�^d@�"O~Qa���y}\ s�� &\�"O��J`��3N�ɠ���1Z� �C"O(	xMR<.���0l��tDJ��""Od)a�L�������	*sB�\��"O�x��W/ƒ�1cȞ�5F}�`O��$f�8T��m rΒ�0�AA�(,D�����X�h�����[)¥�G.(]��)�b�����N
@N)	��\�A���B���%�v<�uiB�y��5��k�-(ZB\�r"O8('��V%2���g�1H����"O`����(��P�7f��cMb|3"O�𳫈+$�p�
����N��)��|��)��1R��"s� �=��b�F�VF��D.�	0�6x�Š��`�N��$�(B�ɕoS)����v�Z���hc�B��BH(�F]�xjp�����.C䉅��XDn��:����"$%�B�I49x�H᪐8�"Hz�$*�~C�IE|��Z�AU�B��8�D��5�h�OL�l'?��l=;�b�t����w�İh�����R|X�0���~���a�	�M�����@������pJ.�1'U�q�݇�r�uY��bh�#7%��D��������p�»#��\k��5L�=��!�X��#`�`ÔJ�p ��;�T���GA�}�S��$_ �'�ў�|��N�;)h�A���'v}j�y�`�]�	d���O��\���\��<�JD	Ƿc��<�*O�=Y+O�i+�]+K<��I�k*.��e�'�a~��M�U�LU"��υ3'��������yR3LX���g�,2��B�yBeG�cXꀨ�n)�u�ŕ��yrg��:4<D��P�:M&b�y��[#��U��C,c�H2������'�azR	Nmr����cy��(�l����>)�OnlS
ڿ]� g+Ғ1p���3"O��j��Fu~�5�+W�ns
�q�"O�\aU(O[���٧O�T��"O��y DY�G*&)�%��e�2 �`�|B�)�Ӕe�� ���("W��+�o�4!OC䉺O24 ����`i�ɲN��Op��hO`�	� �j\P3o�f���F�Y��B�	�oޜ��c�P$T�#@��$B�I1^�PQj�; ���ŧ�	FB�I;Q�tEڇ-�#qM�|��`�B�C�I�V�$����}��Xc�����C�	�2�轺�A�~l̑��ZjC�	>�F��r�[�e�r��r�M-��?����B�T�� Ң9�v�x�F�(!��ّ�z��&L�}�Q���h5!��3y1�Q���hf�8 �`,!�ΡZ�lᓢa��D���v!�Č�	2ZA�g��S��P�n��B	!�$�]Ӟir�˙H4�R�.��'�!�D�"{L$̳3cQ6N)��4�ƚH��O��=���}1ܑc���*��Q'���p�!�ă?-F��P������M7^�ў؆��$`
q$�)��i1D�HC�	� H�<�VO�-���7u��B�	
Qx�e5iґ=������G6t��B�)� �EI6\�p�	8eQ6��%� "O��i��z?��1� j���"O�������Z@t"]#v>���"O�M6L :O���4��,j��x�"O�1
v+[+udM1��(4�"O�\���ݚC&��"��u�T"O4x �D�*"�����K٨�7"O� �s�A< (��6�I� bdL�"O:9;'I )��<`ѡ��b�p��"O��KSǑ4#qj�iTA
�x�"O�,�<Q�t��� �[	�!�"O��ae!��DrX��A���@�JA#&"O�1jV� �Fu�S�*��M�"O�䳧`�����S5/�<�r0"O�u�@f �T"5%��Zx"O"q��������*�?�xa"O��ƣK�b�^U�"���挭@5"O.I�W�A���3���-u2�9"O�|鐥�-F�
�2J�("�ҳ"O.u9vd�r/8X�h�0m��Z�"OT��� �s�B�C5�JQ|<��"Oh��v����ÁZϸ9�a1D���bǜ�q�M �k���7H1D�`��l�
vTPA���c�.9��;D���H��i�$`��	U"�H��,D��i���&p~đ�!�F�G�ð�0D�p�M0i�6�г+�-Z�,��&�,D�؁�d��c�@����p� �t�,D������%� �PЧ@o����� D�,;�,�B8��X����e)�k0D���b-��a�K ?Eh�jci2D��CFIT�e� �bA��ߞa�	/D��@^r�$�!�ߩ]�N��n�zj!��M�Y,�t�%レG�f�1��U��!�d�aLy�a��yq,��`+ �E�!���v���U�w�Ҹ��O�J!���i���q�H���L�B�!���X�4R�>�������bq!��5s5���Di/nn\ܣEk[,VY!��?�~��D&
/j�Z�cC �!�DÛQX>�J��`&9�B�9�!�K8�lt+憃��hr!HL�!�d;����a��!�Z�!0M�Q!��w�F�z��;u����A� 6!�\!c�Y��<
��ȳ�B�wE!�ĭz),��T.�)*2eR`NZp.!���2/D�e���%��l���ΧH!�M
�<
�m@�g����70�!��xi:|�s�Q�,�,��#�2`�!���7�XH�����h�aBT��!���b����"R=F�Ht9���&k�!�$L:�e��D��9#���u�!���pIy����y��F�@�!�d+9�F�i'���u ���	�|!�^=�l�f��Jbh���^!�d�G�f�%��Xn�b�(Y!��?(�����Z3i�%��!ۚ@T!��E� �|��uf�2T�^h"�i�oL!��L�*�[&�ַN����0	�h>!� M,�,�DG�CT�UL�`\!�F�V�&��QN��\<����U62O!򤊋^�.-��J^ r&�A��m)!�E78�&d�U-��^��Xx�K�j�!��
F������?
Y��#�Q�!�� v|s���Z�:�!  vf	8�"OUcf�R�]��@�!u��"O.l�p̃�_�Ta2����
�H�r�"Oҡ���X
 -fL8�)4RR$�a�"O�I@geY�>X�B)�3R0q� "O��a$�ͥE$����^Sl(3�"O�����,QS���M� v7�M�"O��i��_�W��#b��(t�"O��r�B�y�R��l�3�b媱"O28�mY�
$�3ՄY���b�"O�HIEi�R3@��.��@��"O�HH��H՞ W�D�"O(�;�"O&l�G���@d��,F'(��	A�"Od��V�̰q˴��&
G	�4Q""Oд�vN^�mR�ږ��(���"O�)P��/����`�҂]Q�"O 1�f��9��\��f��z"OR������)H`i�D��^d�Q�C"O.��֛���j�d�;E��G"O�+�!��'��`����4���6"OP�St#�)e4̴j���z,�{4"O��RB���;R��끁F3ڝI�"O��)����\c������	B"Ox�e��V�BcGjD'(�Q�g"O܁��A�6>���٥�% <ٱg"O�-�f��d;�E[�'B1m �Ȩ�"O����@�2�,���eG��@�"O�BbVq��1� Z\6%"O�h%�ÍB�d�z��ۼE�D<[P"Oĩy���vN��D��B�f= �"O�0RrH�$%�	q�B<�L�9"O&�k�E�"�0HS�F�`�\�u"Oؙ����έK "�g���{�"O�����V��5����?@w �i�"O6E�K��pN\�� #*�85
1"O���B��\���.��e>����"O ��苨O�0ԇJ�% qC"O,��a�mkBU�g�#8����"Of�@�'�ojF(a�]0Ot�0�"O6`H2HD�G���Ԯ��q ��"O�P:& K�{�R]a�OD"Y�><��"Oځ�5F	Kd�Pp/O�L�TL)�"O���gEI>�((���z\��"O@��썵K�(�tϒ�%��01F"O��s��/��ŋTę�y⁁�"O4Њ@鈦"�.���"��	N%b"O�����Y�jhnUzр5p	�a"O��c���5>`�	@ ֜W�f�PR"Oi�Ο���t����!����"O� �JD6�<aQ�R>0�^`��"O&H	׸>m��2g��;��;%"O� � ��@�=���6x�6<�w"O�����0P�ek��P�^�vĈ�"O�J�<oJ$��wMįD����"Ot��  9.7@��)^!锑��"OXDZ k=x����ŇS#4�;"O�I{�FМ( �yW�7�li�"O.��R��TZ8�g���.���"OzpK�$?�����F"g	mH�"OZ���&Ҕ.`9�Ub�0.W�]i"O�� �	ûb��ˑ!ؾ)A��z"O��kֈK�e�����mC2"O���瓕/b���%̶F
D���"O��VK�?!P�qBs˘(i�郆"O�  �"���D$���Z!}j�djC"OܔR�L?� 0���_M�b@"O�l��\eҩ�&��N��Ҁ"O`�y�Ǉ�C
� �d��25��"Oёrcѿ�r`*�ݣ�Q;�"O=���[!Q���36�� \쁔"O,�٦��<�^wF��\$ �"O6��O$|T����O3#�:��`"OfT�0��%X��� ��ޑ&��h`p"O.��1@��,��I����GCh��"O�UY�H�0����bA�R*J���"O�����(;V@:�Cȏ~$P��"Ol��)��
����`��<��e"O:d�Cّ&����-НcfL0�"Op5@@cN�LZ����K܂=8�s�"O��;6B&W4b�A�:B}�"O|��f�#q��[C�L6P �@"O���U7t����D[DT�BS"O~I��[oJ�*��;nh9 "O��{�iS��T)3B�>[�,��"O�� ��N&�t�u��v�=�b"O�-	 �K;U�F���1��ٗ"O$a� A)0#��[�oY�3���"O��h���c���ծ=g��|J�"O�����I������
Q���Q�"Oh*�,����	t̿�( H�"O�4�2�N-.Y�EVr�`��"O�y��L���Ѣ�%A3}ƶQs"O�ܠP�B}Ȅ��D�v��"Oڈ�1#�#����`��<+�"Ox��%Cݩq���B�W�HN���"O�I���)w2���	Z� H�P�"Ol�H�Iđ%�8��F��DE��q�"O�u9�/ؘj�HV��#D�2W%!��V�������+��d[W#˪,8!��X~Z:��	�7�pYZ��׾N5!�M�O^����Y�O�Vd	�˸
?!�䒋_p���䇾3����e'�TN!���9�f]���M�z��$�d��x_!�DF,{��}h&���A�y8����Y!�צqJnH�B��ʪ���*�6�!�DL�����$]�&�(Q�T"cr!���* (Y؇kƕ*X>�+��2!��`Yt�J2V)Y�!3�g\�!�Dp�2�iS�U�V�<H���ȓfa��Xu�R30�ʐ�3�ş|�l��8���ؠ!�/<��j�OD�����"8DPh�*�
R����׀��%�ȓ��(���|d"�!��R�5V��ȓ�����T{�Ɲ�p�O�:�هȓ ������A�I�%�Ł(.�m�ȓ]������V�QJ�Y�fO]<E�ȓR�.��D�!Q�̈���9W��a��`sX)�e�C6^R,±,��8=����	���(��ˬN��Qw�8H�����]q�#��8Z���.VP�E�ȓ&�B%���\?8��sg#�$U�@ ��2.��r�IJ�m�~�z�h�&]�B��ذLi�.���2fL�9+,�C�I	k� ���Q�4	�vQR��C�I����$��.W�Ɂ�#ƾC�Iy-­k�.�7��$1ӊ͏lO����T�q��ԥ*����)��r�^צ����՜!.4���� �MqH3D�� �!zR,�5$��\!$�,{��t��'������.)��D�l]V� ��\�f-�ȓ&���!m@�&�5P�х�5	��S�
a�~���)r���^�h<� F�l�$$PjH�l,h���ɘ�H��	'0����1+�?f���#�ќq��C䉱?[R��4�]v�:�5/��F��C�e���r6@�Q�j�e� kN��d�1��jX�İ�����H8Ʈ@#=R����j��棛�w	�Pn��t�=�������S�;�H�V�ߟ���qn��yRIA>�.�b�l©[1�x�'�W��yª�|����@h�l9��>�y��U�l������b1z��E��y�Eɳ�x c��˘g�,RB��'ў���ѐg�=7��)�2	�5biKv"OI���P�"�P�S�i�.�H<����I�R���s��6t����w�4*w!��J�!46=��� |D�5B���5eBqO���$�
MI��bD��?��0��3B�y��xR�Oഩ/S�<ׂ\£N�p����"O�q�_�H����Q:[-���"O���'���ѩ#
Ԑq����ύp�<���αf#,�#��Ҳ����e�r��0=9��:��M�ӃL�xp�T�&iCY�<aP�]=H��qB�§�͂���\�<Q��=k�~ڃ��"ss�}�S�]�<	�OLE|q�c� g�%J�o�n�'��y�擊>�� -ܯ!��z3͖5�y�&�gy�}���D�	7��c����~��'�f�����%Q�� �,$�Щ	���1��K�ӌ{Y�4J����z���Z��B�	�eq%BI�1yb�e<�B�I&5��D�BQ� ˆ$ҴX�}!���~�t���+A�6�s-/G��O��hO�B�����'�����S"͝�t!򄘚H�~y���_�Sd��
<f!��D>3�:93f�$o?0����[EJ!�U�J�>�c �M�12�4����55��]�i��}��e�_�<��D¬"�`B�	/,��B��@w�t�wlK��t��$WZ��;�����jA��`�i��*A�1�ȓA���r� ��/�A鴮�/PL%�����ɂN�j�'�D$[ӈ�)��97-P�<:��
�'����SŘ�v�CA�d��dJ�'A�,ݶT�#"�+P�|8�F��|y(C�	�T"ny��Ϫ4)fLz�cL9�B�Ip*�T��
�	]�Ī��uW&B�'P,�0�c���"MQ�%[2��#<щ��?�5G�+p&��DJ�1:��&�<D��0a�=���K]4b��6�6D�dX��ϕj���1A�@
�EH��>��������BQ�Dd+�$�U_���c؟0� ��#����kC��Q�,�����<�eeu�(�h��A��-�c�4g+ =�å�OB���C����t���
fis'cΟ�T�>�'�7�'.��ƍ���h�5Wf@����\qbS���|K�KÒp��Dx��)j�LȒL����#�;A���H�K�H�<�al�:v#�������jsةH�*�|�<qAN�0F�	K	�%�A��d+T�$xC+ �~L�*΂!!� �A(9|O�b��r2�E,�V����%z�h Ph#D���V�$�;�e�|s�� g�;��L���g�? �,8���rwR4��յLD��pw"Ol�ӂ�ƖP�<\��e���68'�>(O�����Y�PR���t��Ycg�Ȳ@(uH�>D���-ߑHЄ�ر�z]Z��3%b�8Cቇz� ���Z�47BЮ�J
����'k��).�����:c'^�6g�M �O(��$�:jhX�S!���$蘖Ȍ�&�O�㟰�����17�=��S#c8%2,	!��K�ެ7)��~�b�	t'�)��O���'�)�ɋ-e>�ib��Ǝ$��B�Y��!�D���};C@Wh�Na*��_�!� q�D :�Ȁo�Ȁ��V�z�!��Q�t�ư��ܑ0#v�Y�L�{���Xx�����)|��b �=4��U�/!�O�ʓA�|� �$-(x�ra\,.YJ<�ȓAN��"��ܻw`z�#g��.�p��ȓ	�(�A��we
�ͅ�Zs(�͓��?a2	2-���3��J�_��ٵ�E٦1G{���i�ƕ�`��_�M��`�+���X���6��h�z�G��7R,���r ���?ѧH�)2T���'��w[���R`�<Y�%fs2�B�Bw.��qF�a�<ɂ��"?�J@���'Ny�Ec��~R�i���)���I�X6NU����&G	�n�x��/�O�ʓe�n�Xq�3	s���fW
0>��m���t�?�g��?1G�޻<ج���סY��4[�<y1O��,��P�љYp@9A�V�<���2v�T�e����HçI
HX�ܐ&\�d� Ȟ�d3����J�f�$��7��<�S�B���
P�N#(9�LA���r���=����T��D\<�`�U/rs��r�F���'�z����q��i��-7�xᓢ��(�M�3;}��O?�|&�pK�b�ڒ��Y4�|�Q�*\Oxb�4"&�JAn갹�Ɵ�,�����&D���CFAe���4��t�Be D�����s��ź��д90V� �1D��+hl�@�y�L�??���`C0D��0�A�%d�^u#!��
�x��4D���R%�%��e/	�h��D��!����	3�!;`��T_�y@�d�%a#!�$/`~A��h��3F���c�n"!�D��tF8�37�4,���a�0!�D�8N4	1� �` ����_��!��A/sO*�����p|\�C���K�!�ԇ5�&Q�%��'5�P� W���!���d��m�qD�9���J�[�!�$@�=�l�Q�kL�wf<<"�I�#�!�D�h���樕tv��Tg@�@�!�D���І\g�,�!�c!��r�l�bEH�T�> 0��R!�dȬ{��s���q�.�F˝5n!��+1C��`&�Bz�.8;ď�7Y!��05j9��j��[�Z��V쎹O!��?5Ԛ�h�+���U���f/!�D�a�lq����Pw��"�؅h!�d�*e`�B���~f8Y`7n�u�!�DX�RΨL��7,뚐�tπ7 �!�Ϗ" �������Y�g�9�!�92�:DJ�j�d��1�7	�L�!�d�Hڤ b�E�+	��4j�
� i�!�Ӿf��
7��('#�k$DE�!�D�,����%�&#�ek���5n!��2Ch�U`2�Y�B@�
:S!��ݴ�>H�Wcߘ�D#u���!�� Z������.��P���@tL��"O����jU�,�3f��2>�
�"O��h����T�M�""��jb8:�"O�Dc��^6�	"����c��$��"O��Х@֋l6 ���5{Bh-�"O�TsAgY
p0I�Ϗq֦Д"OX�r�G�0928�5o j�fX(#"O�d�7�ʠ,�UӦC, ��T �"O���ܦVQ�h5Cŗ%p~A[�"Oܘ�W�(.P�h($#�SYV�H�"O���g���$�tȆ�͟D�,x�"OZ=c��;*Jh�� �7;�*D"Ox�k�*�/\Mb#F6��X�"Or%pqΙ4�#�Νm% ���'���b�@tѴ�*�H�0�9�s#֘���J�'3z��7H�z�q��Y�=�R��'!ꥣ��(~��Bn��OO,8��'���SaH�,\�rM)>����'���R�L�5�V$��J3"�u��'�xMo��V��);7@�*M ��c!"O�h�m�)4�j���;G���"O@�Cte��'L"�bvN�2�䁥"O�h�fMG�Y�F�y�Æb�P
�"OD�:��dc�p���ʁE��p S"O�|� O�]�8L²�\�}�z<��"O�T"A�
�f�Y��ץ<�H��"OJ�:�!j�XDR��PRj�#�"O��I@�X<�䭳X�/L��"Ol���+���Te�$v4l���"O�jt쏙z��e��
��n`�Y�"Ol(1��H#��R�G��R v��"OX`д�]�b����S,r��\["O�����M�B��a#���f��2"O����P��q*fHV�_=p!3�"OjA2 �%�>Q	��s���"O�ts3�G<g6�PgM��#�~�R"OXt���-e%#q�ep��f"O�}	����-���5O	�c4"O6!H �ݭl-HHT�N�l
�|��"O-�E��0.E !"�^1J�
ۧ"Od5���ٽP�y)0�X+t�X=[�"O��RT�ڋ&T@PR�Ό$��<�C"OF1j��Э3pzQ��NH�|���D"O���u��@\!t�J�PR�J"O�[£P K�4��tm�;�l��"O*eI3��W�������4db��"O��@��1O�#��B�J�4`R5"O����HR=6R���%�@�tJ0"O�eS�c�:��e��ǖ8���-�y�䆓"dq�堞:*28��a*�yR$��n�8�B�B�.*4�����/�y�&}�Q��%�'Lc�<�fN��yBNߨF�����u�CM)�y��& :Y+��90�Xv��y"��s���ӫ��~-RVHV��y�×
b9��	�H͚}�l���U��yB�:�d��ҫ�.g(es�
��y�O�L
�ג&���"�(�y��F�|�V�s�*�6��|���3�y�"M$�!y$��W���EC��y"fF4E΅2sdJXQF�ѷ����y"C�'�I���"W$p�*"(�y����`�D���Ʌ�Hʔ!����y�LS�#���Q��T�A�f�*�K�-�y
� �%RF�)�t��'�!S�^��"O�<��A�<�Vd�F�#a��<3�"O���R�&'F��`Ƃ������"O U��H�V���pe�!h�l\;S"O
�Aޅ�|��
O25B��"O�)H���+�`���k�)�""O��'듒,S���W �l^ ��"O|@$����1��	LO�( "O>��!��+U|l!�q�V,��B"O�q�F�q�*�J$�,`�y�F"Op�Ԯ�+`k�3%�L���"OXȁ�O����)��
B�z��v"O�qb�����7L��ڞ� "O�LfCw1H���E�d�z�"O���'b��S�
�׃rh��
E"O�Mc��G��QIe�Q�wn��G"O�d���
y���0�V�d�V��"O2� ���$�
1Сۋ7���Ä"O�����w�r�!@]u� ò"OL�*���mP<�� \:+�PA�"O��{�{#d�`�bĊ0���"Oz�Sqʞ"�>�B" ��q�4�SB"O�(��#�!:�����������P�>���]�0���?�X���0ܼݫ oٶ:�hCR�5D�0*#NԪ}G@��R�V�yf�A�$Pc�	�xb�i�d0�3��\�(�r�*q~\�{F�D�V��ę{JPU�� -��XYS)��޺��$��'0B�x��7����Ĉ�	�0���%���xP�X���BPkܐ(q
�m�3O0ɑI~Z�<j����N|RܡB�4D��*�Mf�!��a�l��I!&�/`�� �^9x���b��?ك�2_ě����\<���y5^Р��գ�y�ߪF�|�#D�)v0B���P��z��=G~��R'�S"R��@)� �+E�t�'�D9��GT�(����rYZ���n�;&Vv�9�[����pR� �V�8}��ڲ"�7P�Ҵ�q�F���×!I-.-�tM�(S��S����c��hN�Z��J����,��ct����&!<Ĵ��06��Or�Ƞ�@��j�}Q@_�H�X#�'�TM[����M��	<~�6��/J�I�T�!T�]�&����W�=M����d�D�A���`L(�!p�ni�D�>m�nXPŅ�-1;2�� O��<�l���"O��R�c��6h,�Y (�n����Hn�~�RF9�A&��v���UjF�)`��'�-�ݏF��-[�&� !V�����#{�Y��ɞ( %���Y�C�������	v�`�SBB�`I !�R@	o>�\Ƞg�?".��Ox$����'�\�a�Ē=ehJx�rCc�]���D�I�ңj'~�����I\9�fQq���"h�$�(��"2��Ċ2v�i˥F8�0=ɱ �"H��p�V��bX�U�HT:	 ��)N�l2�d֥�<��h��bLK;��r��� E����d��D2��$�l�9�'���jE�P�[�!])z�R��4�Ra9�H�vO4�#E/���0�;P���~���x�V�'Gj,�
�� �u��M��C�9/ڐ��	6y�h��&n�4����*;ֈ��I�8,�W�_�A���3�H�0� M�j�5�'�3}ҁ/@�J�P�H�ES���$�фҸ'_TQ����(Cv"J��D�q��j6×�7��H��C�)s�)gɟ�e;h�*�/���>a�D��}=��
��e � ��̃N
l�Wc�*C���I&@�=�,�O��r��<�<��'�Rj珌�>�$�X�L�uߪ�
�'�\���+����d�>��m˄]�T�����+
L���+ڤ��'��i��W���t��qCD�0��2Q+������<9��F3R,�ɐ!b�wL� '��5;�YѵN�I���T�[`�y�S�8}�	�!���v��L�B['\xPc�ײCS�� ����CP�����)V��dxf�7%�p!3L~2f�%=֢��%ťFLN�b��@rp��m�]FT����n��yss�Cg�P�ƙ�ad:x��J�1+.����h�06V>��@�oX�yvP�`q�H�_��[e�M?8K���5�,4��@L2ZA �C�@Qh�丸�bH��<�dA=3�����[(�h�H>��KO
Y-�`ͧ����B5�~��3�E����	�4�t�����C��3P��-E�A��
�i�Tn=\$�2/�IK��s�I)�dW0��%����LYF��B��@�D����2�S*�r:�CP��t�	K�Z,��u�� ��TY]D���d
4uC�I,� H̠�)޽=:�0 ��AI�ٓ�\���;q�R=xt��A?@؈�^=��	)?�Ҁ�*0F�9#�G�~x��g��]8���&L���qP��l��k�b�L!s��҄=�td��O6>�<9�0r>m�C�G,b�x"�K�	`�x��;B'>�!#���	t�^Tp�B�-7>�	>� ��0F��\bh��mn�,Y�"zkN��un�?�M��
O��3#��v��X!�Vs�H�@bǏ�1 ��t��!��}a�q�Nۚ�?90ΗD��݁`zu0�o=rH�i�F��A��C��0
�L���k_�x:4�6L��(���IfI�=��]�׃@�h�P�I�e�X��c+�z8�gy��
���X3�f�*DH$� �p<�B�M&J�q�@a1?Q�U�G&pZ��'E�"@�3V��$��Al�`J����<�c�G0%'�ԡ��נS?��97`^Q�dU���ݞw�%��"�jƺ>��3���`����-��Y�5;�o�3f��
�'�X%�)�:o�vXr��.�[�(�2��9_ C��*f8�rv�(Xv�}ޱC+�	�Rh��Z�c�N@S�`'$��GI^�	��`���6=�����b���!�`�
��I�+% �#d�Ӝ��gy2(C6"����W5�4Ճ`�C���<����4�6OhIQs~B���Ϗ=6��G�7��0�����a|A�|a��[�5w���:`nY��p=)gmݷ3� �s���x��]a4.L�\ɜ�bG�ر]��:'�G�Ɛx���>]�1 c�A)�%����8��'���c�}��dy� �A�q��T�"�.)�F5s��:n�\�"O�Y����0��K�G�L���Cܴ�U)�(�0Gx���Ծi`p"}�'K����JV�m���`��\w��a	�'Č��ᄩhn���A�U�ܝ�C�0@�����Jy 5ݨ�0<!ǄR� �8�DD�m��a
�p���#�l�$~�Vhkv�L�L�iK%��P�+�L:q��	�I�!�¼p�X�;��E�^-���@�/�I�J69j���a�L��o�*S���4�c�'�����w�j`� �;]�X��8E*	(��:k�~���D]:?��pӓD�e���J8OԹ��H�v�/4z��c�O�E�r��o�h����%���:��'���2fM
�-H�|Ir$�gg�	���$"�'@�YR�Ͱ5Ί!3ц�&&��Ĉ-x��
�!	6ԍ���^N�Q�0��'��e�� sA\�7�M��H�.�qӗlf]~�`�<���*Y6|�!�D_�>ε��A*{_�a�'B�[���E�TJ雲�Ҽ2l����؞�PDX�`�}ܧ~����ՂP768L}�U@�,��̅�)�f�Z5�\.=xِ`�(E��d�R�(W�����a�;�*�+�W��C�tO�� hm���7��%	*8;��M����� 	�t��VB�5�b�uP�7����i"~p@�jF�Y�a|�ӿU 8i�eb�j��$�U�ւ��O<�k��$\,2`�f�-��V�jk@$���TY̪��F돮t
!�O1/�L+
0eBj���J�DJ8ZW�5`�КfnF�S�O�P�2S�^�w�P7L(iR����'[�z,�5%�	d��c���z��>&H^�E��M�՞��}"
фu�"XaQ*ʗ4�$	�U�]���?1JQ�t�8�x���(ZNv\�UE�1V����Ƀ�x"oҏ���b4`����ؓn��y� "��sd���i�@�C��%�yRDB/\�p L���d�2�M7�y"�֊,�� ��S2ʞ(�H�y+ǜO���"fC�$�hV�D	�y�)�l"t��P�J�
�f�B�7�y��I�^1x����^2n�Å/A�y2��u<��d�C����å@F��yb��	*����)K $I��� �y�`I��TcR��5���A���y�Ȱ-
��Vb�+�\Z���;�y���R	9f��%�8�4a��y"/���g�6��`��ES�y�y�.q����!����y��M��q�'l��|��h��OT��y��5:��M)1N�D;r�����y��[�@x�H9lwD�	&�yr���9�Uae���
�*\��j� �y"�E���*��@w�|*�:�y
� 2�c�:,�҃㋗�\�r"Odr� �9̤�fh!wFE�"O0���=��S�G�)}P)��"O��@D�?�*�3�I�	�)��"O�	੏� �TX�&�;��U�"O�A#T&��zW��QK
C���%"Ot�9�*�8�N�aS
�%kh�"O�1����z��Xg	��*�,L�"Oب0��10T�Jg���6"O,�S���S �Y�%��"��i�t"O����J^�la!?p�РR"O����j�}|а�6�s�<@"O��rc�ɜ!�*d��G��z8"O4M����[3�U�' ����p"O��sA�XL����P�W`~р�"OF��p틀A���Go�p��8g"Of��1+�JCt���Y8=袍�E"O4؁��Ll�4�v>d�;6"OZ�׆X+l����L9�'"OQ�v� 3������~���"O��pC�����7����"OԄ�P�.g<�`��Z^�pH�"O�d�ŊXP���T���=����"O,|;Ac�q�i��bK>�*�g"O����㏷||�p�!�2c�r"O ���A�>?��qvCN�z��tK�"O�h92�d��d�!_t@L�!"O��;�G*0t���B�Au���U"O�XU�Ur�j2G�]@\)��"O 1�qj�-x�h�H10!6�"Op���M]�y��8q&DR,��!"O��'j4�ZbD�#D���"O��C�ֶ&t�e��l�T<�"O��e�L�.��]�&)�~�Q1�"O��M�=$v�{�ʕ4��x�"OB��m�#
����T)2�|p��"O|i��!�X��qʏ�/��Y�"O��* -��a�Ȅ� ��*F���D"Oe��M9-±�e���n��8KU"OHX�򥉃x��p�3���rQ"O��9��-Q���[���sTI��"O��TJVN���2CO�0�Ե "O��R�KE4�>�C��T� M��"O0����Xpӡ�v��AX`"O�����݁�N��%@�b��Ё�"O8)��N4o}���$ݑ?w��)�"O$�qL�L�dl�c�rVx�`"O��r&@�%_���p�hM�`�5"O�ڣ�C6 FLPW�[	cO��c"O����b�䄸�� ڐ5b�i"O����*�ms
��	�>�N��"O0����"~=.�k�	0^�mpU"O����"L<��ς�U7�@��"O���w͕7o�9 �N�#�ظg"O �w��� �����G�Z)f�*�"O����lq:.lc$��47���@"OxU`T���l��(��H�o%���"O(=	D,�4S��X�+�3$%�d2�"Ol8��`Ǿ`�v��Ζ� ��"O��Z3�.50��t�@!2%�A��"Oڈ�Q
R4K���c��/4iC"O� �T��A���P�O	�2nh�7"O^y��̌�6=0(Sv��3C
� �"O�D�Dn٫YK��b��4�P%�y
� &���Rl�>��䅹,P0�"O�$z�O�s������O���["O`��q(	m0<��P+��l��"O�l�4(�y�fxᡇ!k�^��"O���C�Sc���7�;p���p"O��fŒ�9ʕ��F����P0"OJL�cǣ?�V�9�d�>D���k"O�0��ىXr��sŃ��!���p�"O��@%IW�n�0C��A�'@;"O�a#���!���!MIdk$@a�"O$��E��a4������@"O�	�g׺l:��C���7"Ot�4
���&Զ?Ӯ`�A"O��BRK��b+�h�j��O����"O�гD��2X�, �KƼ$O,�7"O���)�/s���ԅ��d���"O~��ej��%b�����]
~lm�P"O�T���G�V����j�[ `�""OH�7+Ξ	lH�#��7?V�f"O��r���&�Zt�
�w)|A�"Otr�!V7ɔ�S�'^�A�y�3"OZ��I'p}��g�LG� 0"O�-+�(�.g�*�@���<>:���"O�����W����se
����`"O�E����o��ɇ)��Z#"O<uB&/ sܕ��(N��dU B"Oֱ�#�)���a��(rڑq2�>��j�P"���?}9GH�#p'�0��d�� *D�0���Y&!&��d�ЫF�n!�oWc�G�d5�T/7�3�45V��a�$�(p�,�p-�2}Z6���B�M��a���=st����7��udW�>�xPD��0;
^��$��m�� CɋE����eEV ?�����I���)��2�{M|��
׵OA>��rCP$�}���t�<�E�Y�5��H'�LR�����Z���� _v�ؤ!�aĈ?��E�*��]�i�j7-E0L%~��5�Y��zgC��ks!��;:��b�3D�P�Jg �d�c���-QT䨅�q
��gF�=��*H>��w88`�.�)WܮU�!Й�4`���'��p�)n40�)@��:Cc̦H),��į�jGȩBta�)03�x���>Y�HB���?��E ,,vɂ�U�i�tJSlO��Ol���+
�[P8�¥�@�w�z�j%r���P��]��lҌhg�<S��O앺��[�b�jT+ӓ5c�j���	O�������pC�͢0����0D��?PLy *JA�'+��U�aȄ)D�F�g�`�Q�ϻb��i(�!���y��F�Z�`�نdK�L᥈�? ��v���L��,�.� ��WD�W+��qA�>�O��N�RD޿_��ɉ�$�CN� �$|Op���ȁh�N<����3J�>]�BM�]v}�!�AnV��NS'(&̜1�%7}2I]g��?��f.V��aeLÓs4ajQ�
B�',�Li`��+_���C
����O7P�ʧ��q6^�q)�'PJ�@��'�h��QJ��O�4����g�&��򤅏*-�@�i�q.x�+�)MP���b@�6�D�)���@
5�Li#g B�e�$H-��@ "��A#�>�z��t&=D�HZ��RBr�9d�w�$sՀ9�H&��-A�
�3KN�,�bj��X��I3V�i{DPD���H�@��Ç�FT�R%�zF��+歗�t��Z�#�;s }D�_�a�~�X���l?� H�����>�'��ٲ�.L�M�v����-y²9��'
��PM��X��lh�AK��2)��/߰�ȅ�IFX� ��/���l����%ݚa�&�;<O�x�Wh�#הuخO��'l����O#a��"O^Ac�A 2^(�����\��ɳ��|�nƭY�����H�t�OȦ���a�h�KĝG�ͳ�'W�u����E)��9�ꉋa"Y������'�4X����>YшW 2�yx��4��F��}h<f�AX�ہ���xe�ͺ:e�Q�a��ռ��d��u0�`����`���=P�y��^��n��V�^}}bH�>��JBhR�u�R�r���y��t!�A8$'�s1�����'0� �j�i[�?� (iQ��
0΄C�hB�5��9�w"O���"o�):���/"�n�8F���/�qOV3��Y��겁�p3^pP�ťrQ����/��'rdA�V��>�5ҫnt���G��
�r�YRdHH<�Ԋ\%1;D��G`;KP �dL�J��A:�Ä�p?WD��-bhm�@ݼ>HPq� f8����؃v��4Qe����3c��.�u2g�J�o"��� 4D�|[c��$��b��2xl]�&C!}��zo���B�B�g�Ъ2]?�y��5m�ʡ����<�#3D���!cñM�،���k�t�Z�ǒ�72�'����%&�'0f������y'�wh�� Q�n�T�XV���Px��I:h`����8�V�����*}��`1G*x)r��O$�9���W�X�R���� !���*�قC��0��
5��x� �c
<�B�@d~��0s�r���Y$l6���4 �.>`��m��U��9(����?֊�BĥS'' ��O���ʥKFrK<K�H��(�'4>p��m������N�@;���'A��@	�9yԉ�Ҏ=^�$�t��
���$y��	�iI��H9�`��Lr�����e�>������ ���u�1$�������Bh� ��'�:m��_�f!�`d����	?t�V0�����gy��Ԓ(e,K�lM;i���1#���<A�,�;k�ObcD�i�X���9$�`�R*�0D��0�� Za|� � ��2T"�Y�����Q'�p=�!�ė)m�[��5  ��ĉ�~LeYnފV��`����x�CC9�J,�*B�
���CgO���'��I��N?��� W�	q��LSE��ɜ��#*� l�&��"O��� "Ļ�d���6j�D媒�ެ'H�ː��
s�6u���iTV#}�'8�iZBS�L��3
P*���Z�'~�%����"y�lL�s��QP	�ڢ:�5��*F</l������0<qR
��M&lI6gTU��`���r���95E�,2̀�ҌH*Z��a���4b �!�Nʊ	��8P��I�!�Dڍ6��Ȗ�_*xǫ!��"ZXz���ܮG����e����EJ�'1Mx���)�����1[�Ytv݅�pb1X�D�J�
�r��F3@�$Rw� �T(�A.@:l(+d��c��Z�z�@�O�-��a�>[Q�JU��v����'b��yƌO�`kTq@��Ͻ9����4+QD�0Ɔ����W#�)��d�rŔO����B��<t�W
ܖ˘�hă&�_� t���x��MI̘�C4d���+B�0m�PCd�H�7O|˖ ��Z"��(�(��Ķ8΀�`+�1��$b��$�F�]}(��Ať��� ⛃b�@�������#��}%��`�h���^�yڎ����p"��gL���1mKd\�����&`,QYFdYܮ�yN?Q��̈r�7�Z5�֣gP^������*���	�x �#�%x���
2sO�|�J��6:t����(;�Ej�̒�h���d��4��5
~LD}��N-��A��L��LA�OTh4I5ЌI��heP��QZ�'�p �#!C
_P�#�O�[\��'V��'ܠ{z���Z��}��$Q2��à � 3g�� E K^�<�UAV[rI����7߼��@���Izk�m3Q�����g�6B&ҲC�&RP`��,st=����7@"ҁꝃ���G�����+���=��v%���񄕂}�Јç�@ ��8�ȓF%��Q6��	P���{��_�ObZ%�ȓ.O���Թp���k3b�����ȓ.	����&�� Q3
s�=��r8jq�B��<5<j�(��C0;ⶵ��% 4��f,��#	'DȈl�0�ȓ�q�@�A�S�$�;2X@��?��|���X C��ن(�bl�|�ȓV0��
�ܭP�ְq��_"��ȓ[b��,�D� )�cK�k�܆ȓ	pX�`GNߐ� �(�j۸ن��	�F��`f��l�o�L�h
�'�B�A )V-����b��i��!�'�Lt���F����@f�m��'`P�0@S��6E�t�݀].�!�
��� ����eҷ*	P�"��^�P͐�"ORq82L�<F�Hx���U���z�"ON隂lR:3�ic�P�3�t�@"O�a�ě�,��pp��@�kz��%"O��{���B�\21f4x�1[�"O�e��BʎzB�R��Ǟd����`"OZ�*�RӚ�h��?9ݪ���"OP����
ZBr|CK".�@���"OFA���R|��)�]�k��m�"O杈Ҭ�DAvp�3`E�s�\9)"O��j���y�މA�*I�X��p"O����}��s��8�p\��"O�(r�H��Mb�j�![� �"O�xO4{�.����"���@
�'<��������U�:y��j�'bC��}�<�s�45�T]b�'j@A`]::G���3bڑ ;^4��'�q�UD��g��xC燡l�R
�'�dq�S��9l��W����	�'-��(���#(�
	(�eG/V����'�t�k㌔.�9æ�$V����'�Xl��܂q��U����C�����EWf�:6�%M��H@$��<��0x�-ؠ� ��ȓ2�b�17,��s$`�B���5�Ќ��q����{d�i�y��4�ȓ*�*	9W	׺z$x�&�	M�n,��C�D F�O�P��m���
��P��d�l�j0��92��BJ^<W2P��x8��&�ЫP���Z���f�B;|�'D��Ă(Tt�S�O� �:��C����K [�0�Ҁ���a�f�b> J?c �eF����ߩz�pD�V�1���qf��M����Oq�����T��D8�e��i�`\��
}
3b#�����+�n3�%���k��F�8�M�5r.�{��@~2��=o�L�çy�A�$�5Y����jˇ"�*D�'�Z	�G ՗A�E��'p|��s�Қ��#�a�*H=t4�E� �	�: ��槈��� �ɐk�|�2��Y�+8���,&���HG/!��)�ZA�P	��4Ӫx!�@Ҟ�cv(��hjs-�<Y��`>����e����YF������Ym��TQ+����S�'|I�k��Z �p��C57�|��'�7�\�����ц_j��i�V�?��O�l���]�|�t��b.P 6J܀N֝lZ������M+�FC�t�S*L|�UG�
T[�Y�W�]�:k�u�Zq��`��yӂ���0�ư(�$��JФ��}rBQ��'�]���
v���Ib��'��8yj���O\�b��ɇ��BD�Y>���$n҄!�7-Q�R�@ �G�T��]�������S�O�`�r"E�{ڀ� C7)@"�c6D��1�%(X��pq�;e�`L@�4D��"/��z�H�	!?E�4�Z�?D�<:��=b���`�3�*�)�c)D�X"��    ��   �  4  u  %  ?)  ^4  �?  �J  �U  �`  l  �w  ��  �  W�  �  ��  ��  ʴ  �  V�  ��  ��  [�  ��  r�  ��  k�  �  h�  � � 7 � � M" �( <2 �; "B aK �T �Y  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9��CZ���1.*��5���#D�������=9js����]>+-B�I�L,����ơT� *S"0G��B�I�<w<̉@���R��Xrȕ(Uv�B�	�n�t�hՈ7Cn���ӳ;�B�	x�Ψ3�E�V�B�ʑ�ޕ-bB�	�K��� L0B��h�'��O�`B�I~����b��L�5��£~�B�	�0�dq�  -Nz����� 9�0C�0>a1%
�y�N���.M7@B剖+($�w������Ο&|`!򤂰V�dS�D�
��PZv�I!��"���㰁L5=�����	�!�ӄA��a Q�&�ʀp`�0#&!�$\(�����N*�Z1�f��+%!�D�J�ݨ�H�UwP5hd�	!�$C0�d��#��1a��ɷ*���!�$J�gÔ�[��,;�2	:D��J�!�d�c�\���HOOj��q��o�!�R 5rZ@
T�� ]VH�RbY��!�dI�{g)#��MF�EQ�J�7_%!��= G4i�� �<+������5�!�D
�[�T��"D�*��Mr�N�2w!�$�aFڈ�&�ذM�t�D��l�!��.a��To��6�F|��,	�v�!�DQk�m�D"��W���wN@h�!�X��1R�/߽`v�S!/Ìk!���/uӦ&�(__�Ո!�ǖE1tܙ�I�X�Ļ��̓�!�ԉT���k�E[*E������6#�!�d�zr��h!ꖰg;l\��cT�t!���k~�X oF>@����c�#�!�8H�Lk��7�Fxk��R/�!��Z�^l2��^ a���Rf�L�,�!�$�� .!���"S$�*�.��2�!��0BYڨp� �:8P���KȝW�!�*@�X�Oފ?g��ॠ_�)�!�$�P��+D����z�� E�!��  �!�O�M ��#Y��"�8#"O<��"��5Jf<a�AmJ-�Xt	U"O0�8��+��k�삓���"O����HM6��JB1[��ЫD"O \�!�Ðq����g)B�6 �@J2"O��FG�`:�}�C�F#f,�3"O
��'ME:,�qq��s�(Eg"O���	�;y�t:�ɂ��)"Ov� 7�	+N�H ���K��� "O��c�F�T�ʁ�Ҽ'�Rx�"O�t�䃋1��xI���VfRYj�"O��KU�_�(>���!މ�t�b"Of���m�3��P�N(8���a"O�J�K;kм�2R�I�Uh�@#"O����_�QbKZ 2�pq�"�-�y"#������O�sd	���J�<�SN��M�غ&Q���9Í�y�<�Ed�GW
�f�[A'V�vd�\�<�㧗�E�����8��3&U�<��M�*%(0(�Vː�@3��Ӥ�v�<A�C�{c2(HW���>I(�)v�<I�_p� �S7�эF$�4�4m�t�<�6�Ì�8 �%�{�$@Fiu�<����6D� ���υM)	��p�<YOB<u�N�yt�@&t��(0��T�<ag'\�*�%�fW�:�Y�fmEl�<1��2�(a��N�9�"}`�
�p�<����Z����(�^�m�S��G�<-����bA�E�� ���_o�:B�	H�΅���b��y &�*|B�Ig��X#�'cz�`DO؛t?B��1V{����ʑ*O$� *(�B��#)b΅1���:X�Q�/P�3NC�@�j1r�ԈS&�mSG�=X�C�I x$�A9�2?\����όv�B�I�o����7�ю Kt��GB��"aC䉇+J�;���:~$ *�C��S��B�	��0�3vӤ2�*!� �)��B�ɫx8�l�tB����Ԛ��p�B�	�VV�IP�MK�?�@rFY.!�B��;2?��rq��:��4�6!ҵh��B�	�s��*�F�30z���/Q2k�B�I�M�l�8��	)���q�[�B�ɽy�Zp�L�	p_�4y�$��]@B�	�B��
������r)]�~R�C�I�O�FT��K����RU�Z�͚C�I0#̓ �¥ 
P�qW�T�G��B�	�M��{�E �jlDp9u�ǵ��B�I�CJ��Q%�Գ�bH:ņ@�?JB�	.?_$���ǉ@�~%:��Ql� B��PY)�r�A� "���iܽa�C䉻>�iQ�-�Y��b2�[Y?&B�	�9���ʄ'6"�����	B剓KhZDJ�"�+H���$�F�FO!��v[\9 �&Q��t��$�̺H!��9b�+������$��
5!򤘊bE:@yb�+��r%�U5!�dX3m��t��^#�̤[��O�!�$��\�J͐�J́*~�{�$F8,�!��$�0'����(0�ڻP�!�dȠ�H�ʋ��(��
�!�	*��4A؊k�$�"Y�^"!��Ime�!���\j�r<�5�Y�<�!�$;MM湈@W�1ʦ��nI�G�!�� p��ˉ�	>R��t�	,J�p�B"O�9IU \�`6� ���Э��"O��kNk]�9���97��8PU"O�E@f$��bk���fF��t��8�"O2T�.� ������Ρ7���YU�'t��'���'��'���'���'zİ�r)�7B�*�����) ��'�2�'b��'>��'���'�2�'��R�i�F���*��ġK�T:0�'��'G��'��'���'���'��QJc�L���:C�T�OB��s�'9��'o��'p��'"�'E��'7��0%i��:t<� ���J��y��'���'���'{��'��'b�'�U��Ƅ[hj��d�,"�u@C�'pR�'���'CR�'~�'��'~���G+�()�a�5���,(n�X�'�B�'��'f��'R�'"��'�v�R�Q0A>�k�U>OA~��'�2�'*B�'���'(r�'K"�'�lu(����[i¥�TB�)������'wB�'���'�"�'�2�'��'y��AR˃(@�����_�}5 ���'���'��'���'�r�'?��'�@���HJ�V�f����O�]0(�'�'�"�'�R�'�r�'���':��'���w�Q����&Q�-7hT�P�'H��'q"�'B��'���'=��'F�i�Dێ
_$x���ַ��Uy��'k"�'���'+��'�2�vӔ���OR�9^��		��=:~V���[y2�'��)�3?y�i �MBŨL<u���Y�I��'��	�T�?�.O��d�Z�������+-���)���i���$�O�ph�h�J����j�H�Osxk�&��qB����훸:ad=C�y��'`��Z�Oz�8���G�z:�偰[;<���#�>Y/OV��.�ȟ�]�K�`�y�i�6�^���d��?*�E��ϟ<ϓ����x7My�x��ѲY�vp����(�X<[`�j��J����s�����'"�Y"��z`8� (Y��Þ'#�I`�I���O"�(A�0B���P+��ĤD�,�O�ʓ�?I��yrR���NE B����`,�j	е�B�+?��o�f �ťT�'o�d���?A�lY9_�t�*#�#��!�����<)�S��ycE���\�J!��œ�5�4U	�_G�Iy��'��O�[XS�H��4`0��C��
`G�$�O.���O�q2V�yӺ���4!��bMQ��VF�!���Dd؊fL[��䓀���dZ�@��IA��!9{yY��]�I��D�O��$�OZ�?��$��\�D�e��f8/Y�%a�	7�M�%�i�O1�lX�AlO-�$\IRF�&��AIb�w6��*1�<1eV�=��İ�䓆�H�:1�m�wf�=W3�,�s��#&a|B`�>9��prFcT�s��iP�F�9A������?)�"\�(H�4Q
��!|�NM�O��~O|]����*�;S�A4a��6-h�p��3`�*�P�O��Ж'��4�w�D�R�.(C�X%;'f�a2���'���Ud��(����*^�}��C�r�'��͸>�O�ҝ|"��|�P|�4��;nи��)G�jO6�lZ��M�'� h�ܴ����	�~t�`� C,8�!`H�.��R����?!0�#�$�<�����+gKʟuc,}�`�O���'�B�'orP>����@�s����|H@�[�%8?	/O���O��IU�'h�� 1욁d"������ mN�P�F��	8ى޴]�i>8��O��O��p�̍t���;��`��X�Od8nZ�f7b��vj�0z��@�x��Iʟ�	ğ��?Y(O�0oڰHvJ���ʍ�}�QjT,CJ��ܴ\����$Nƛ֚���T����j�nyOA��$a���>F���A�e�y"\��	џ�������	�p�OLDp�V�"'�j���!A�JP��@�>��?���䧮?�Ӽ3�*��z�`1� ��y�gS��i!��O��O��E1��f3Oʔ!׆3�\��e�W@��2O��5���?Y�(��<1���?A�陛*�2Y���_�]�>I	��؂�?Y��?)���$�a}r�'��'�bA���;X���k��K�4����$�<Iֱi�7-WB�62=��ACL��,��9 Em�*3��	֟<ɲBY�'��2C�ty��Oט��I�G�r/�?)unѨPN�`����՘h�2�'���'.���X� T�p\���ʝE��U�q����lK�O����O���:�i�Q�T�'�D�ڑ凣A��Rv��y�4}:���g�r� Si���D?���������3	�F��T͋κ���6~��O`ʓ�?���?����?����Uqv�		�:I�T�ݪ.��Y(O���'^r�'���d�'c�"�jZ�W�D[�E�Jm�`�W�0�	ȟ�%�b>	KT��7m��D_�NH���L w�	spF>?��#�F!����<����D��lB~��E�B'	A���o��G����O��O��4���5�I���s�V�!�l�4�F@���g���In����$�O��$�O~Ȇ��B��rB	P㚥p��A��7�6?a�B��	$�S��� ��jcI��m���2��݆Kg,,�g3O��D�O��D�O����O��?�s`��)h����G^=~z��C������ß���O��O2��6��0;f�� EJ�Lx�����## �O���O�� �Bm�6�.?� ��M��x���#h�>���V�@���d��On9�N>�,O���OV�$�O�t�p�ȓq�^�CP��9��͑ĉ�O&�Ġ<�S�@�	�� ��y�d�|z���A�Pĉ��d�����<Y��?�K>ͧ�?q5E���IIREV�sB�CiG�tS�:
Q�4Up�'���,��:d�|�N��}�J<���6����K�"��'��'����[��ܴ_;�����LV����K���$̓�?���?��T�|���ڌ�G�%�%�����p���� �&�����?Q��2 B�)RO~�'A�C0��iD.�HQ',�yT���Ο���ß�����O�xd����_,RX ��y�@��>y���?�����<!�Ӽ+��O�k#���txc!+���?������|���?��49l�<I4��/�LxH@�Ȑ>��m˦���<�H�U��d�6����4���D-0$0�cFN�1���k�-,|�D�O����O<� ���p��̟T�!S�I���5$0����Pd����O��9��Nw�~UP���")�\� 	�/����?pR��G� T>c>݊��'^>��	�Z�ኤw�$ەH
>�D8���' ��'���'X�>��	.[=��U	�(��["M(<����	���d�<�����yg��1`�U��G�=��ܻ�
���y�{�Dlo�&�M%��Mc�'R�L�+���S1.��ʵ-KO��Y��I3'.b��s�|�S���	�����؟d�IߟlpI	��=�jK�B��ȈJy�Ȧ>q���?����'�?�0�J�|C.	q��\.0#��c@����OD�� ��O<��O;�-��CU�7��-��"܇bV���]�T��[�`X� v�"�l��ay2��1έ�PkҧY�𸓂X�Z�'���'��O/�	*����ON� VKKNAu�!,M�k��r��O��$0�ITy��z�Ƽ�	Ȧa��e´A��I����i��X��#����o�[~B�C�<�lL�S�0u�O�g�I{J� Q� �fH1��Գ�y��'-�'���'c���R�w���Gxf�8���Z!eW&�d�Of�$�q}�Ox2�':�'��I�4��fjnŀ��H�5�
���-=���O��O�Qմi>��7t�.}hg�y�={�+u����w��j�q�IEyr�'O��'2�.�<LЄq�5���q�~p鱣ɕq�r�'6�I���d�On���Ob�'*E8��W�z���X�&_�NB�`�'��Iߟ����S�t&F�JE�"uҠ��zAWReb̫�J,P %Z�[���*�2hEm�	��৪�p b�	�i�	ȟh��ӟ$�)�[y"Go�,)S���XX��	-bMļH�6OF��?�RT��A޴P�.aX n1�Hp;���P��
��'��F��W.����< ��Xj+���jyR����[��/en�$��h]:�y"P������Iɟh�	ҟ��Oޒ�*�M?M�L0�������)�>����?����'�?9�Ӽ{�I��
��l �b,A8��ʦ��V�ORO1����#iu�*�	�X�1�W;�,y
���7�@�?Yx٩C�'C�Y'�̕'��'&`�1�#�d���Hl�^�2t�'{��'��Y��@�OD��O�d>Bq���.Q8��70t�㟌�'�:6�B� &�X�Ď�$O�x!�-�:DQA3?�Bh]�J�v���%��N�b����?q�9�^�U¤j�R�åE!�?9���?��?َ���O-�JW5Nk][AHT.{�f�S��O�u�'�"�'���4�`�ˣg]9ZXڂA�
���1OV���O���Qo?87�.?�f8hŲ�i��	c� �h)���$шb�D�H>	)O���OP��O��D�O�5 � 6���&R�ח���m}�'���'��y��#8�Dp�C�È20lb �շw��	��@�	F�)�>����=Hf�؅��+�4lY�Y!�|�V�w�{��f��O�ʓ�F�C��N=l�J(�(D������?i���?!��|�/O!�'&���B���F���j�^�թ����'"�O�˓�?����?�a��s����:F���M8H+v�4�y��'��7#��?M#�Of����% ��O$-*����� �C>O����O��d�Or���OZ�?]�!-�@�(��TL�4g�M
���ğ��	ȟ� �O��͟�$����.Ó{v�%��1��u:Ԩ	X�	�t�i>�XPaʦ��'c��0��6b_��c2�M�<S���f#�J�Xy�����d�O��$�O���O�:������	�#] 	�%ڿx����O��I���ڟ��	�P�Orp٣'L����2��;[TdX�O˓�?����S��EOH�{'.Cs�r�˂�U-v]āAq�1uқ�n�<ͧX���l�k�"�HsC �te�i��Iuр(�� ��ڟ��)�STy�s�86վV$n
����&q�<���?����?9��T�p�I�`#h����7`1�=��G&t�	�|�N���a�'�&��1-X�?餟� ��	c���v�l8�] #5��S5O��?����?A���?I�����ɹglД(�h�kpF%@�/°/O��'�r�'"��d�'
�wv���,��dKr��#im���ia�'m2�|�O���'�|%�i#�V�}lj
1�#7���*�Fܙk?�֡
�<8R��7iƓO>��|
��vdjE/?6یȩE.V�a�I��?���?�/O���'���'r,�6����+�BAzn����O�˓�?����ᖽ�I���'{8&\r��@~�"��O���Xֵi^��~5��'&�ؓ�(QeH�M��}i� @�ko��'���'"�Sߟ���
�6�z�����/�<�	��Zݟt �Ot���O��$#�i�����߬��E��(��v�s�Ds���Iϟ�̓1<4mZ�<���>����j�?���I&����j#x�����s�Icy��'���'��'��H��X����Dj\|�S(�1_�	����O��d�O"�����E0,nݐ�G��h�%�/",j��?����ŞFTz�p����
:�H�ẻ+��9
�����M��Q���$��=���"���<��C�l<Zt�5�Z�
Q�WD?�?)��?����?�'��Vt}��'�P�c�]H��ّ���&�P�П'q"�D�<Y��?!����I�.Ҳ$��|�1����Č�����M+�Ol\�2N��ڌ���w�b���(�8B���b=!����'�2�'hR�'�"\�b>���S6��Qf숌Gi���w�����Iݟ�9�O�	�O��.����5V��X' <@<$u���X.c��Od���O��1l6M&?q��%�-Ɋ��0���ڎm ���O��`I>)*O�i�OF���O����D]+bX]�S'�>c� |�t��Or��<rQ����矨��@�4ju�Ì�7�ع��	�Lt�'u�I��͓��S�t��1Dw|	�,
-3�.=S����z��CdK�X���Bs]��S�xB�w�	-(�9�'k��� 37nԒ?���Iϟh�����)��fybc�Ё�F��$*Np���DܲC�-�t?O��d�O���1�Izy��'��"jZ	:xy�A L�T,��	�7O�7��uz6�4?%�����iG*���_���-p`V/,��HK���<����?	���?i��?!*��X�Q'��)Oȩ`ч�Sx���G}b�'�"�'~���4�80Q�:`oh����˷$�T�9P�KӦK�4[����O�\y9�i��ėARX̹bOC�iq���'k� �Ŝf�
��x�`�Oʓ�?���U �%KU �<N�Q�QM�H�,<���?A��?-O@5�'u"�'�b�U"��l����sd��1VjY#s1�O|˓�?����|�hh՚M L����:!� Y��?��\�{����4l�I�?�[t�O�d[mW�Q�ai�y�(���␅S"��Or���O��$=�'�?e�L<i	D�c�'B6��$:#���?�T���Iٟ��	d�Ӽ#ЈƕtJ�9d�Q�;�����<I���?���RO���ٴ�����B���F����ND�sC�f覀�t%�����d�O����O�d�O���Z��D�[��͘���z� ��PQ��+�Iş�Iʟ�%?�	;g���kV[~\�I��
%>��ܗ']h7M�ڟ�%�b>y�2���cyPy���}��Y�膈Q���:fǔuybfE�8L�IS��';�Ƀ6�B��FPu·$�FÈ�I����	����i>!�'�`듅?s� S�����ٌ;m����Cҫ�?����'��ɍ�M���'���b�%y�"�_?.�i��SS�d�s�i��D�O�xJgꆉ�rD*�<�����ӅT*#�|�P�TpULt�r(Γ�?y��?����?���O�^��!� +�Hϔ^qN��p�'���'�d��|B���?YN>�恋#V���SW�t����a�l�'��z&�Р�M��O�y0��B	5J�m3��O:$�!c�Nt�>� ��O8ʓ�?9���?I��p����,T$"�^�������q��?i+O���'2��'�BP>qs�+��Q�;�oݸ!�}8��-?�.O�o/�?	M<�OH��ƒ)S�LLg��	7��epv��.p����vN�i>!��'S�%��[�lQ�d�8��B$X�y$�Dꇢ��T��˟��I�b>q�'�7Z�.͒Ÿ�a��h��l��B�u���Ot���Ov⟰�'�7���R�@e
���z���ĠWE�m��M[�-�;�M�'�BjS�U�d��S&��I�I��,�W��e��s��^6X�(�Ry��'���'S�'��^>�B�� �N�a�G�;�Ɖ�3����d�OF���O��N�$�O��F=]+ ���	]� Yѭ�%yM���Oj�O��O2��B�d��7mh�0ZAl��z���#G	�qm�1`c%d�L��Jݸr��� �D�<!��?��E�Q�XX�-N�0�pv�X�?���?�����D�h}��'��'	*0�S��LWl\(� �x֠QZ����<����?YH>��Ǌ2:TıVNŢm����ǯ��<Y��M��,���6�MeU�h�Ӂ5l���O� ��Η3������ �z��O���Ox�$�O��}2��)��z��B�u>�89rkM�E�)�b���П ��̟4�?ͻ`���DK#i*x� t���.3"L̓�?���?1�ڟ�M��Oݡ�&����� :|�1bPr��u���'$ �mK�"�ģ<���?!���?���?Q��^�5>��Y��r�&@���$Pl}��'��'���y�Y�c36 `�bW�~ �hS��]�E��	3�M��'퉧�O�L= E`�!�ɀۧo�e���L�7A�!bpQ�$p%�	0Vr��G�Iy⃕�Cb4!2O#h�֠A�U�2*��'�b�'��Os�	���d�Of��Ě�0�,�s7��:�dP%��O��$2��vy�'
R�'��X˳�;`�X�B�-`�� �-ՙ(���7O��E7�2A��Oh�I�?1�]p����!lY�{����Ҫ^�.�	ߟ������ܟ���`��DR��V9f@a��[�����?�4$�i>������%��o[M�h��&ȃ�h��I`��ӟ,�	������=��?T-ֶ1H6u�񢆕�ࠈ� x�`Ͳ�䳟P$�ܕ'B�'�"�'J�(YƭA��D5S F�$D���'�b_��Q�O���O��d�|���61#jAQU�� ~��P(b~[�d�����%��'�1�I�#M�6%�Fm��Z	����7x��޴C��i>ᑀ�O��O��k6CT�L��2ti�)�Պ��O.�D�Of�$�O1�ʓ���f 5`8��j3n<nulES�Ȅ��y�S���	c���$`��#5o	�Txb���X�I�|9Q������nzK8�9n�p~��V<�h��'f���>N��P��ā,b�0ف�.V1����Uyr�'���'
B�'*2_>R��W)s� �KR��$q���!�0����O����O ������O�H-��Z�dݩh����\
n'��mڄ�?)M<�'�*��!v5hݴ�y��]	>����C9^Z�4���yn Qr4���0!��'s�I�d�ITi�i�Fj�х�r4����F�˟���̟���Zy�n�>-�Ms���?Q&@��ƈ�T'ѩ]5��+�/����'���ןX�In�5�֭Ц`؊t������G�.���9jp'���M� ����Nq?�����X �&(��Qe,H7_`��S���?���?����h��D^�J|Y�%���w�V�1��N�
���$�G}��'u��'��O�.=rrg��+_�p�H���z�$�O��$RΦ��Næ�͓�?ѕc�R|��ɝT詪g�J�.��pp�-6���M>)(O@�d�O��d�O����O�!S���;Q��f�W u�>ܣ.�<��\�l�������t��� ʱ�c&��Q��7	*t!�fyr�'?�0��iE!?{E��'K�����3w��)w�X�K�˓�h�����O:y�O>�.O,]�����+�I"���e�����O4��O����O�	�<yAR�H�	6[%d��Pe�8)֘zW!	H_b��ܟ��?A+O�o��?��4=Ҵh����#r�<��" _�^¶9��{�ٴ�y��'���9'�?�y�^�,����Yh�B8Ǭ�4�ύEś��g����ڟ@�	����I���K�q�]�4)[�w������K�?)��?A5X����(�Ik�	6
w�xruK͒\��,bV�	O8`�H<Yּi$"6���3Ă`���	h��DL�iԪt��
�1\߼�{Ql\�8&����'�p8'���'�2�'�"�'�0U:�ӁSP>%2��l7�����'z�P��٬O�ʓ�?�)���:�[�f�b�A���WfB(PG����'�6m��q{O<�OL�	`E3+�B�@�&(��HÅD��x���+�ca�i>%��h�;cj�'�ٲq�E&t��4��Ӟ!����' b�'d2���OS�I-�MQ&Уa��Xg�\�k� ��e���<.O���6��vy2�'��@��E�4"�zqgዐ�Y��'jb�T�pG��0O��䊘sD^���'$���fQb�ʒ%W+\0H�I���gB���ly�'��'���'o�S>�:�d­gz���l�kU|�[`k�����O����Ov����O�N����t�Ⱥ�Ђf��X2����O��O1����r�x�I�Xְe��e3h �]�p�,�^�	�Yn��F�'�P�%�����'�|��� @�d�āhU$���"���'��']"Z�TA�O��d�OJ��	�:]�u���N��'��0�⟘�'�R�'��'��t��Ɲ�6��R��)q�	Ø'A�Q�,_�A� �2���?Y��'�,��ɣ.{��b�b΍qqb�c !�;q&L�I⟬����8��i�O���Z����������,��0@�����>���?�����yW瀸G���2��׀�$@`�ֱ�y�$l���	Ħ�;'o@Ȧ�'� `�@�?�{�i��ª�1�-ˠr���)M ��'�	�T�I�8������V�����k��I�Ь�����'Q���?a���?�H~z�tZ�9�˚(J����K�Z��*�O����O�O�O��s��+	\^T�a-	�W� X��M��<)@��@U���"��t��CW��ty¦	VD �BG����T�K:r�'<b�'9�O�	=���O��Î]&U�qACD�Bu��>O��0��yy��n��q�	�12����*�$ �%�6ݐ@.܌y�6�n�F~RC��p����ӣ
��O�w��k荫BIz�ٓ����y��'�b�'s�'v2��9�8ڴ�'\�X�P��_���d�O��D�]}ʟ���=��Z�}�"��B
�+�:xфE�֨�$�|�	Ο��E8w
6�=?�#Xu�? �p��ӴT�.ȇ͗5V��r�̊�?��3���<���?i���?)�$ĿUJ<���C�3(\,i�Y-�?�����a}r�'[r�'L��<�1����&�дg��v�`����������S�����6�����;3`� ʴA�h�(h���*�`�C�V��ө:��MX�I$v�Z�G�X�b;�댙q�A�I�d�	�p�)��dyr `�T��0��c%��c���zI����5O���?ɋ�X�(s�4[t�0�EJ�<&�&0���V�<Ųb�'��V�A�E�6���2�G^�x���NyR�M)n$�M�"&�zI��fR(�yR�@��˟��ٟP��՟|�O9��`G%՜i>h` e�z��9��>����?�����'�?	�Ӽ�� ����+S���j�����Ku��\$�b>��)Hɦ�̓d�U#����KF�k>���pd� �g�؋F���o��Jy��'��Ŋ�*F�3�ٍ]�*�[׎ Sn�'���'�剐����O��D�O�P���˔z=��0�^#F�^���-�	m~"�'��V�1�D�Nv`�Xv�d��w�9V�x�J�O���!/�X�L��u<�i^��?�ub�O���jA�B�n�J���,B��iJ��O���O���O��}�;E<1p���)㘀� %���\ 0�Ga��ş��I�0�?�;`'H���a��D�p�ׇG7~���?y�4��F
?�M��O8T*�!�
��X�����(��z��IȒO�˓�?����?���?���EsΥ����9elR��[�F&P�P-Ob��'������V������ �P��=�Ă[*����O���2��)H�jh��R�ª4�b쐆'J�E{�Iu�V|�'P�,�a�j?�H>�(O`Q�(�}^	(���:�M��g�O����O*�$�O�<�BS�����XΜ��#�ti�ٳ�m_����	����?9/Ol�$�O��Ą�4���H�
ʤa̒P�FD1Ѯ��g�p�@�DD�q��?a%?��� ZG��ڕh�'�r���	!<]���4�	ԟX��ȟ���o��}�s&�ÊP���
T�S~+��b���?i��g��i>-���'�t0$f����Aٵ�n�%RN�G�	ʟ��i>�1���æI�'��!�,B��ѓ��
r'�`u�^�1��"��'p�'�Oq��'l��' �];�J*i8e�e��U �,���'lR�'A�dӖ���OD�$�O��'��XnO�i0� ]!�"�3�'��6m�O�䟄mZ���)�|���v��(!ş�iG�����1K�Xe�"�tȚud�-����  ��&���OZ��d�
�+D>� D �`T��O�O���O����O1��˓7 ����v���s�� �l��x�ƥ�y�[���Ie����$�ǦyZ#��3����v G�W�<C/�?�?1۴޺���4��ĖU�@qk�'i�˓�������\BuP��ʍQ�"����d�Oj���O����Oz���|���P�X�
#D�A&� �5�H:"��؟����$?�I���J� %�P��&����m��uj�a�ܴ���!�4��������hӘ�Ij�!��
�oV����	������'�fI'�ؔ'���'ĺ�م�� �V�Q�BL� 3��'J�'�^� ��O0��?d��Q�NX�uO�=üJw����'��8�M�g�iy�OJj2�V�5IȜ��1�����S� ���LbD/�k�8�/�|�"�F�7:�L����h��Jן �I����	��D���'3Lx ���R���+�H�F1��'����?���?��w��"��62���F	j�hd�'��7�D���A޴O��q��4���2_�����'VBq�$�	�4� i�s/ݫj@���0���<)��?���?A��?�0)dΐ����A�S3b��k҅��$�]}�'1B�'��O0��5Q��x�ͮ��ē��D�	��M�i��O1��ly��ʒ�/��D-�̡W�L*Q����7 �n��I�33D�2��'i��'���'4�:1FܿY7�#��P�I	��jv�'�'����S�xk�O���)��2�I�x:=2�L#K�����O<�\�'�r�yW�R=.̈�臆� Iݰ��V���S��Ӣ�i��	F�Nţߟ�������b�̛&���2�uz&Y'��$�O��d�O8�D�O��D$�Ӝ (ܑx`i	�H������;q@"��Iȟ�	*��4�F�d�OD�Ox�`c�U�BIsӍ��E-6�[!(!���O��4�i��xӦ�ޢ�0�fJ'Aܜ���l��+?̵:�;o���W�\y��'x��']" ݻ$?�)�dl�T��h���߅N�'��	6��D�O��D�O&�'*�D��1G��N���jl[(���'��Iʟxn���S�T�ݤi�t(�RG�R���?DQ�%�����.�.�	$^��S%S"&Pz�Ʉ&�c@�d\4��T�J��0��O����O����O1��ʓ(�Fo� a�bH3$�0�,�]���'�z����'��	%�M�w�a_R���M��:+l�ǧǘe���kӾpa�c��	��2O�o��4��|y��S��怪&dL�H�>X�����y�]�P��������`���Oi�5��ge�r��>�By{�b�>9���?����'�?��Ӽ��Ƃ|�0�.��\����bj��n��M}ӈ�'�b>-c�kBϦ��S�? d8JbKI�IA����ힰFrnա5O�TJ߬�?A$�7�d�<����?���߫`�t������W2T1���?1��?A���}��'���'�����Z<ŸiXD`�?V�� �B��<aD�iE��$'�Öy�-s'(�w�j�F��I�I#xgF�2!"A| �@$?���'�d�	'8U��o�lp��
���+��0�	͟@�Iៜ�I@�O&Ro��1�p=����S�(�j�!��(��	�>����?q�����y�ƕ��Z����H2���%����y��uӖl��M�c-	�M��'��]����2�3��O�9[>�C!*�e�R��s�|rZ�Vjӆ�d�O���O��D^�7��2z��V��Y�*�+]��ЩO��$�O�$.�I�O�U"PDԛ:s4��֊�.Z����Ǹ<���y��x�Oc��O�59BA��$��EgNJ$u�ώ�GM�ʠY��ptN��:�R+�d��~yC�5h�5��cK -L��k0;B�'R�'��OE������O�}j���>ʊ4��F���FF�O>��(�	Ay��c�����٢T��jL|{!�����;��ϕ'���ll~2��8>�.���_��O��#lU�1��o��Mv�9�*��yB�'���'���'2�I��H?���#�&�\�{�h_�.���O
��o}�O�"�'l�'��yTh�4@}�{��C�	 ���3�|��'`�OJ� �&�i��	(;/�-��mx��	D��ACrN�j�~�|rW�������Iӟl*���P�r�H��n��l9�����IZy��>!��?1������A!P���
6�U��������wyBgqӜ�m����S��+��L�J��F�ĺ�T�)��貲�LѤ,�^��S�m\�h�y�	'��2'�u�(:�%��kw���	ȟ(����h�)�ny"�`��CD_^<Fɛ��?nC\��3O��D�O���5��Ry"�xӆ�8��a�0ر�
8�j�8�cɦ�@۴%f�<2ٴ���,�:<����~˓O��ܡ����S���V�<te����O����O���O���|�a��rM�a�/��-�����>.���d����$?a�I��]d�.他hȒ|� ����Z$7��TI���ٴ$����d�O�)Z�v4O�u:Fb��U>=�u���/�,�Ɂ-1b��'�f}$��'��'�����J�v��$8�D�O�p5�'�'�"�'��[���O����O2�䜆3���@�-�6;�&h���^M���'!d6-���l$�hd��6�C����ᇅ(?�O��,SX�Q�O���+PL����?�D��" ��G�YV�xQ�	��?q���?���?���9�8g�A�Z��PѢ�QրP�f�O���'w��'T��4�b�j#JE�$��d���_D��t�O��kӈ l�*0Iok~@	"lVl�Q1J�x�L$X�6��өVP��i��|�Y������ �I�(��ğ��U�PB���e�0A�����h�iyb�>����?���'�?Y⁌�P��	��g\|�35�M��$�O��4�4�����O��{'��F��܊�� kO��Y�_.�7�\y��Ίp�pq�������ԧL����+t$(���B?�����O����O��4�
�B;��蟨�6AՀr��U��A_�~����GF�P�Ig�����O�d�OR��"� Mp�����v>� �!_?�6�!?3 �^En�l����{'�ދ/jfR.�/X�ƅc���I��I��\�I۟����.�G�t݈q��#u���]��?I��?i�T�Ė'*R�|r/`MZ[�痥G��	hG�C{�fO(�o1�?�Ӆ��1lZ`~2/>`8�}e��~y^�;��֛s��hH "ğ��|R���	�T��ğ�:��9F��u��i��]rƝ������P��SyRB�>���?�����iƑ�|��6me�H��J�a��	`yR��&��o�)� �t�t��"��O|nU��F�.�ag�S!L��,O���?I�3�D�+�P��h��*m��OE%?���Op���O���ɸ<���i̬p(^�&o����̢,<]`�'��	���?.OΜm�*z��KQ�]
���N�
^�Y���Mf���M#�O���nD�:�j�<��B�O�.�" ��
a``ړgH�<�,O*�D�O����OF���O�ʧh�N8x�S)K@��8�ϢU&�X��Y�L�Iџ���v�'�?ͻ-�60�Tj�T���@����L$�X����?QM>�|2�I��MÞ'�J�:u�C�����L��Б�'F�p;tjx?iN>)-O��D�O\���@�W�`�r���#:U�R��O��$�O�$�<yY� �I����	� �"�j�'�Z��Z���6>(���?.O>���O�O4@��� ~�T�P(W�?. 9�Ж�h�@�?m�s�a,�Ӈ?ia�Ɵ��r��|*4q��L�M�ޙ�@�Hǟ��Iߟ ��埠E���'�t��çØh��u��L�p�v�:q�';���?���?��w����W�7Y�rXf��~'"}��'�7���ܴH6�Xߴ��� >�rH��'\�H @q-��w��1ɑ&h��K`�%�d�<q��?���?!���?�:V ��5�L<����-V7h�ʓ�I����۟�%?����=jD��dO,K������^�;b�'�.7-�ݟ�%�b>�i-� ��yV�L8U�x�"���ݾ��K�b���/�>t�b��O��3K>�*O��F�I�^��@���z��,J���Ot�$�O`���O�i�<��Q�0��61��Z�E��5���d��>ABd�I�,�?�-O�In���?�4;�f�P���O�ti	�D�`v�� ��M��O�u��ϣ�:��2����P��`��0ѺMS +ۑ2���9O����O����Ob��O��?�9V�ML(f!s�Ӧb����'KRڟl�	�lk�O����d'�Hȁ�A�`m`�Ε/L���;�D�ϟ�}��	��@��64?��hn��z�-�
B=����O�$�+�f��4$��'��'�b�'����g�;�V�1d�ªS�7�'4Z�T�Ob���O��d�|:��_�AT�QT�9rT!�B~2Y����� $��'\#*D+��πf��AA1j��=��5�J4r0$�i�4/ �i>ɋa�OR�O�H8��UZ��SG������O���O0���O1�p�Z��ȉr����ɟ h\�ţ	�y�P����O���d�Oʅ�W�ؚh�0�'dP<p�Ҡ���O����Yo6�=?y������I=��Ǉ?n蜙�Ccؕ��g��y�^���Iٟ��������ߟ��O�ܤSv�H� \��#K�w�ԍQ�ɤ>�,Od��:���OD�4�
��2HW&wz`��fa΢ �tAs�Ȧi����Ş
���kܴ�y�I���4�' I�U�l�r�F�>�y*I!{�8�I*gc�'�؟��Ʉ]Ҹ0� JBf:y�5 �'<k�h��Ɵ ����X�'X�듃?����?����*b=Pl;!�\�(P�9p����'U�		�M;6�'R�'>�b�%B�"`�l�ĭ�~$����O�x�b��+�N���&��O�?���OT)�Zo}�`hW�"<m� ��]�?q���?����?��)�O�0�D�1���Ѵ \>`&����Oʤ�'��'�b�4�l�HӌP�-k�`1W�>�n�9O�]l�?�ڴ#� �ٴ���חz�\��'3�´��曧eo"��n�D�j�a�	-��<I��?	���?)��?	�^�t�J�Ň 4� HX�O׾��d]D}��'02�'��O1�
c���#A�0�x�W��,���M��'Չ��O4�p��� �<\�����)F.`��+x<�sQ�� ��6E��G�Ivy�M��1��La`�^�40fO�f���'���'��O��	����O2�F���<�����,[�X��S�O���2�I~yB.v����	����'
<L��J7���&�������7�0?�w��/pe���R"��'���℈\�+�CT)	l$@����<���?y���?a��?����F�%�D�����F��|�U7[j��'@ˤ>�'�?�����	G�ыt�O70����*N�Q>�ْP�xAu�����`5��|��G��cDާocv(�W�޸U]z���͉ +E������䓪��O����O(�䒫m4�,���\���lw��vj��O�˓g�	Ky�'���/���B%�G`�5���_W����女�����S��ˊ�1p���$��3�d)��ۆ9��X��ʃs���@c\���1) ��s�I�,:,�k�Oԋd�0�D3Mgz��I��d�I�\�)��ny�)b�,`B��>���Ó�@Sf��g;Oʓ�?���X�X��s���ML Nv����C�dEh)�	������ئA�'�D�c#��?E��@R2�TY[�AHB#A
v<��34OH��?����?���?����U�.j�=�v�9~J(�bE�@�ק��4�?9���䧓?��Ӽ#�*��/��a0g��k].������?����S�'}����4�y"��8�iQ��&X�B,��K��y���(�}�I k�'*�i>��	�E�R�zv$A)�� ŤP!<3��	���Işx�'���?����?	
�=��h��K�7�N���Q���'��Ɵd��Y��{�6���H�~�Ƽ�cL=?E��^��1���?~�$�|Z�"�O�$��@>9X�/� #a�,��:���?Y��?q��h�h�d��>�i��A%%�R]����U��DKK}��''�']�O�n�:JUQWLU�Ĵ���G����O��D�O�s6�}�0�5m����)���X8��	�,�p����#�>�aR�V����4�����ON���O�����&S��t)`����+e:�����p��矰�*T`�o���`N�pd������D�O
��>��Ɂ,Wr��y���?Y��J��R9e�Y��D��R�ɥr6�ȻB�'��%���'b�$�`��+%ʥ�.��UѺ�q�'�B�'����DX�tʩO���<#��@* h�w��)�.A-^���O4�Е's��''�A[/����HVS��d¡�����T��i���w�X�V�OLq�6�N�[�bDX�O�8	��Ȫ��{��O��$�Or�d�O�d=��s�ƅ ��X������?�2e��ȟ������D�<Y���� }� ��b�9@�A�ܽL�BH>����?ͧn `��4��$@�" 9q7��F^���A�#V�ęj����?�`�%���<ͧ�?	��?�ĠD��$,Q ň>4����"�B��?�����r}��')B�'[�S {��i�+� Lbd��D������O��D:��?� ���a���Сr	��h�G�g� ��/��i>�	�'T�Y'�dI��q5���1д�b
؟��	џx�	�b>�'�7O3s�m�󋒈%����?#9�<�����'��	ΟL%`�4Lh�K)Y�!�Шr2��ğh�	1��n�Y~�M��T�y�		�Z}�q�ABD�߬��5��	��<����?i��?9���?Q*�fA��C�Q�1��+@�-`�	p�(f}��'��'��O���yG��02��0��$Q��������<�X6M��|$�b>i3q���͓S`���uH؎P��s�B*`J8�Z���ص��O6�JN>�-O��D�O��S�� 'mx���[�nܪ���O���O��D�<	@W���	ğ��	
n�\d��	�9?S���R�-R�\��?y-O��l��?�J<YRLݳH�L�#fA6f�l�+���f~�G̠l!.�]���4���C�ӟ����'�2�Ƭ�0�p����Oд�{��'���'\��'��>��		A⎌�Q�I	I��k�aДjT�����D�O����OB��]�o�F�
7&(h��+�p����������u�hE禵�'�����B��?U��=�Dz7���i���'4�I�8�	���	� ��*�z�`0�S�X�E����g�F!�'���?a��?�I~��Lx$��8Bƾ<!�C$uo��(O�o��?iK<�|*�	��H�J�k�B�;9:��Cb�!A�.M PK�����-�0m���R昒O6˓�<�s�Қc��[vD��}�А{��?y���?���|�)O�=�''�3|c�lB��!*ޅ���c�2�'��O���?���Ms� �+az��#� 
bR^��fFU�[��ڴ������ ���l똓���� ������ 	�̐�S�?>���O����O����O:��"���ɼ���	
�%Z7$�e�L9�Iٟ��ɰ��4���d�O��Op����6
��%��[5l	j�ɩ�M�b�B  ��M��Ox��$�w�\��`kγH�mB�#P4�ح	�����O�˓�?����?Q�bX6��)O#'JJ�Ў-Ť����?Y(O04�'?��'�U>�g�_�-ނ9KQGJ?h�RL2��s�(��p~r�'㛆,+�T>��W��%,�Q&CB'8�4 �{O|�Pb�7e78\���T�ȟ����|Rnƒxu0�:'퇮ޘahw���@��'���'C���_���۴`R0��iL$qxu���׹:. ͓�?*O�O�<	2�i���I8*��]C��L1f�����pӸ)mZ]�T�m�p~�M�*��A�0f�剃E*ubփH�b#Y6]�C� �	gy�'���'�R�'dR[>)��C��:�f�P�`*G�=�3�"����OV�d�O���D�Ӽ��
$F ���l
T�� #� ��?a���S�'3`�\�޴�y�D��{ Fȅ�eJŎˁ�y�Ȁ�p�L�������O��d�:��K��/T����+ը^�L�D�O:���O���������������y�(�1��*�n��c�Q�	�<�''�7��ͦ�I<��i�>m�ܛu�X6T�nՊv`�q~r��l�ˤ䀇d�O���Ɇd��R�[o���v�Okp�؀��� _��'cR�'j��Ο�Rb霐-��iHUF�x00d"�����ON��<H>��Ӽ��KL	)��# �}V<�ʔ��<����?���P�`�hش��$�/�!��Ok��a��<�h=�s��;I�Mz �|bZ���	ߟ��I�@�	ПHi$f�Q)�PI�o��q(�)SEybD�>���?����䧏?)b���J0����E����5������O��D7��I�i�F���������E������{c�w�@=�'����n�Z?1H>y/O�4��d�(,˔فTēn��O����Ot���O�ɡ<��W���I���0�v��xR|����%>H(�'oɧ�\���ٴ{%�6�g�v`��]�N6θ���Ӊ	ߔ�;ӮJl*�6'?q¯_����	����'��;R��!�1 �Ofy��_�<���?���?!���?)��4J�*��#��r!ُTҤ������	��4�����O��O���P�^n/�����v�d�ҁ�_K�	�M�d���􄂘�Ms�O���T� "K�7`W�_��h��R�|�~�(��'@v�&���'�b�'�2�'���`�b� N5̡P�m�-&8��t�'pW����O����O����|Z2,��O�@�"��O��@E��_b~�U��۴5��xʟ"����Ѵ "}Qv@&"U`@��k��ě@"Ɨb	���|�C��O�%�N>9�͖���a L�,��㢡^��?Y��?!��?�|"*OJIn��~D��Z�CĈt����(�7Q��	럀�	����?�/O��o� b ��f���D�(�^$J�����tn�K6ZnZl~ ������_'��2w d�� h2q��	"|���	jy��'���'���'D�\>���JS��	�Ոϔ3^�x��E������O����Oʒ�����O�N	�p��"��0S?؀"�˾W��m��?	N<�|څ�X�Mc�'�d����R�����,�P �'��0(�	����|�Y������P��	di��Re�kn��h� Jğ�����d�I]y�>�*O4��ۡt�U�LP2m���a@���hO��8�'J.6M��%�� �$����".�@I�E��6A 5���)B����X�@���ڟ�r��/0�@b#T���!��k����I�@�I��G�d�'��iS֪߫r垽�b��{=ZmK��'�j��?���?y��w��
�$W�1��A���F1p���(�'��'7�րO ~�����,���!r4�$+T�oକ�� 69�6q`W��Q�"A&�|�'���'�2�'C��'*NMH��O;sc�#tl�)T��-��V��X�O\��?)���HE�%��5�'�T/8N�()T�S-�� �Ms�'����OJ{c%ػp�Kp��-�6���I�#󂁫�Q�H�PNN�K���D�	ay2�X�C�x`õ ��+�����¾+��'@��'��O�割����O�� ��]�7��������5�"A�43O��D(�Iyy�gfӢE�Iɦ��l%����aب���j�],@�lb~��Qk6,��(C �Od��1%�����U����%
�y�'�'"�'�r���:B^��q��W����������'���'�듖���O0�O��jG#��nE�[��%�ҩ+��&�<Pݴz��'`0\�޴����k4(q#7X2`R�a�2Wx�`g�S�I�v�Z����*b������@z��:��ԫ+�Y
b��y$@p��$Y�]����
�4]
����߳k2$��gV�[�h�r�&��pR�e�ߐH:H5��.ir�	�g�ԥGj��)� S�O���b�Ň�W�5��d
.)`���nH�7_v�B`ܱZC�����-ꮄ�3�,Z�M�F��8DT�amM�#wr����US' �#�Π$2Ы
%^��吶�] $ ��:5�� B�X	gO�Ub��Ŷ7E�q�R�/J�R �tn�u��a	Wc��\T$#���T�xX�ʒ�KM�����-�?�@�i�2�'[B�'�.��N�3&�L� %E�}$�ѳ;�d�O��|��㟠�'9�^���Ο��	�"+��h�oZ��$���T�ߴ�?����?���n��	�F�AC��1��V�L�?_&qߴ�?i��y���i��䓃�i�\��lU�Lcr�� �-Bj�	�M�����'��'a�,�>	,O�e�f�ܚ
��qnT71x��凚񦱢�E2��򉋯H���O��!E���g�̺�*�&�Aa�����Iٟ���ğ̢�O���?��'���I� �9dt���g���l�"Pێ}�6�y��޼�y��' �'fh(S�ʐP�6��CF�[��%��nwӨ���OX��'��I�<&�֘�T��G
�uČy1��/N���m�^���?a���?J?A�J��*l�U�V�Z�g���W�`�Ф�'�	�,%���I�@���w�@�aH�PG�a����.OV����;�x�	ʟ�I֟�$?M�O����֯��"�0R��ͻBw,X�ߴ���O���?9��?�W/���$�����Ȝ�;h�8Q��YM~�ܟ���ٟ�`J|�EW?��I�}^y㠅	6Xv-X���cG��ٴ�?�O>I��?1��G$��'����e,W�7�Q�C
��SN̦M�I꟨��g�H�	"����O�D�O���Î�O���	��ҝt��0{P�MP��埰�I8[dhi�?i�O~];]	tB��Ŏʫ]�`�شx>]��?a��i9��'8��'�v�xZ,�c.M��½�&��&]�>��G�itb�'?����d�|�O��U9�'T�Y\Z��˄$tS�=j�
bӜ���˦��՟����h�O�ʓ'��cP/B�?� ��M�`/�8�a�i?����|����<q�/�2D���'�%Ƙ��9i�I��M���?y��?��\�L�'Ob�Oܥa$��C� ���e4RL���ğ6m"�dN�X���O��d�O��s.$cx�Q
���30[�<�1�榁��ݟ\c�O�ʓ�?�O>��)��t��m��E�v|���?PBr��'[<욄�'�|�'C��'�~*��B�լ���'݃���7��٦u�O�˓�?�O>I��?)#��+%����ϓ�T�Ź��2F�{�5̓�?9���?�L~�0���ô��"��!a5��A�H��X�P�	�� &�T�����'����U�ݥ4��cՃ�n?�1�jU�y"�'jR�'^�����O_r��^�����åh���;�ȟ�^�6��O֒O���|j����3��UW�ǶD ���;6J`7��O����*N�d�O�t�O��'Zc<<� &\��L�)���4_d�YH<+O��d�O|�����P��F̊p�����㑜M�(���i�$u��'��cp�~���M��?���\hd�:N��Ń4�RW��T2�o}����?a��h�O@�S
��6I �t�JRKS[���LK�k}�	ǟ ������џt���� �t� �ڵa�#Z�4M��	�,.\�'��,���4�ʰZ�������Bf�"���K9��A%`ߙ�M3���?��?1+O��^�� �5M|}�s�G�[}V�Hb��8c�MDx�s�Q�<?����?�;-0�1XOδCǀ�qU�WF�Hn�����IpyBD�~���<®�y�Í72�:)�HX�|�O����	N�	ܟ��i>�x�8]#v yt�r� 0���mZgyb�'0��$�O����4m �N_�Ao`�*c	�C�6�Lr�$p×����֟�[ybПr��"i��Y+��r�jL�ub����i@��'��Ot�ĵ<yB�Ц!RbdǔA���ƃN�K!x��Eʝ�y2�'jB�'�Z����O�rdG4h��;�A�
tr���e�ԋ2;�7��O<�Ot��|������E"����� 7�Z}�)O$6�7��O��$�p6˓��i�O0��Ok� ~M
�g	,i�$�0r�	6s�X�b�xr�'��'B��"<�;_�T��c �kQ�x�s�37�)o�#����ٟ�y޴�?����?9��J����m��̪��Q2]�ba��ؐ`|V7��<���?����T[>�R�d�jѐ��r��c)E>5�a��i��B~�`�d�O���O��'��'EZt�ѓ@%+��r�O��g��DmZΟ0��֟,&���=��b�����5(3�IyCHA�)�R|�úi8��'y2�'|�)�J�x��(	j����N�m?��Q��N��O�$��9n����?1���?i�wa J��w|M��#V"x`z�	��i���'v~O�S]�	>P�F�k?q�N����,?��*J<Y�i�����?���?aI?%"&N�Hވ	�GߵE�X���*{�D&���I��$$�Ԗ�uGL�Dt�)3� 	�<��c�J%�MC��[��%��?����?IJ~�S=�$x�ufU45>nIX�۽lv9�ƺi��⟈�'���'�b`�?���^w��q6�S$%�@��@��Laz���?���?1����'Q���۟�X+����%�ګ9�%�g6J�^6��OB˓�?���?�����<����~ҀD(	$P�sIωg|�RP-�M��?�c��<i��PS�S����I��d��iA�wƂ�5�[��<���$�OX���O�iS4O�ʓ�?	�O{�`Cn�z%DT�2JV����4S�6���?q��i���'���'VX�Ӻ�R�EA޸�n�=n��p�$E�禽��۟��gc|�l����|jƕ޺� �bk�����G=s%P�9�N��E�ɯ�M;��?���?9bS���'�p����j�T���z~����fs��9�7���'��' ��՟�z���+9t��P㐩T7V0rh�2�M;��?9��?�Y���'��O$a�u%��#�2���jN8��"��7!K�d*G-��O����Oz]�$6P��Uꢌ<XTx{�L榡�	Ꟑ��O˓�?�)O��ƞl5�� �ء2&#*y"��Y�i�⬏!�yR���L���'��'����5�AH#FA���f�	/֡��
�M��X�@�'IbV�D�Iڟ ���<u&ӱV���C�d���(e���n���Bg����	ϟ����?�O�6�6P ��T�������..6�<�����$�O����O�ȇ4O����<sz k��=S9~�2!E)G����O"��O�i�;��L}����5��;���0��n]�QI���M{�����O���O�ɛr3O��d�����N�#���q������)s�����O�	��<OJ��@~�t�'�R�'��EX��D�М�#����3ɴ>���?Y�e��Γ�?�)O �(y�iJ#G�^	���i��6�07�P�2���O�`l���<��ܟ@�ɥ�����!��]x�`��A�D �t("�i��'�~�[�'@��<�.�t�IĻ�tpT�`���ұĽ��ۥ�M�����'�b�'y���>y-O0�y6��NY�ID&KM�y��h�٦=c`+?�.O��'K���Χ�?q�E r��њ0F�HTd�q� [�`g���'�'N���>�(O^�D��+���S����MV#@2���"�>�,O�h��9O�Dx�5���$�O�D�;H-����±Kt�l�h�X�oZ՟��	?���<�������Ok�G#�ɣ0 �4lq>E�ׇI�Uz��
.���IA�L���ߟ��I����s���	���r��uT���cB�^��6-{}�U����xy��''��'���&!��E�D��JI�	���yb��+1U2�'s2�'��TU>%;�O:��Ja�T<,f2��FA�,Y6ms�4���O@˓�?����?���w}�`ÙE�� ���aT����ʚ0�������	ן0�L|B \?���E?&-��*�������4L��4�?�.O��d�OV�6w�i>7-�S�hS��Z4!"��b�MJD�f�'8«[,�y��'N��'�?i���?��.�0K�Li�#�"��A�A6<�	����ȟ���O3��4�"!��<���c�i�PJܩ�M�ӫ�<!��f�F�'}��'DR��>��yX��aRE�\��g�h̒�m�ן���#[����|�e���+��އ-"5�P���B�f�{��V¦=�I�M����?����?)�T�̖'�>�jч]
&<@���.,n�	���`�R�7O���<�+�.*r:����� P�	��Q��i���N#R� ylZ������P�	�����<����~�+�� 0tL�m��\��ՒT�����D�<�B��<I��Y�|b��?Y��[81�T�
U&l
QhJ�{B\ҵi���'�들�d�O���?�1.8�L+�B@\X=���a���'�p܃�'8�� ��'xB�'�b��yZw�<(�r,��V5@�{s��m,��4y_�I}yb�'��	�������l` ɒ"[?$ŀB�B�(; ��s����,.���������4%?� �O��X0��n���b]͔a�޴��d�O���?���?�0���<!���#3OƠ�`F�TgX��s+�y�����?����?i`����~*��3Oz��f��,w�HT��+)Sb�궳i��T�L�	���I�վ�IT�ܴc�-93&B�$3���a"P<hz�lZ����.²�	���A��f��O����a/Hy���6a� �$F�R�]�'�"�'0��/�y]>�b�7��mO�U��k�<H T����릡Cv�(�	=�M���?	��?aP]�֝5�����ע*��M�C�
U07-�O���VD�Df��'��Ӻ3�*ם_�ڡ�U5!������~��6��Or�n�������I���<q�� H쑣��I�
h�1O.2S~-���i�a�'<RV�ĕO��;�O�F��QmjP�)T���0�M]7��O0���Oz�a}Y�p��|?��H�9E�Q�c�2��Q��@Uڦ)�	��l�� am��I?uh�ڟd�	��8�FC;���{r�Z6u*r5�Ɲ�Mc���?	�^���'�"S���i�mH�̚�=^��R�?�8*��>��e��<�3����?I��?y����Ӻ��f43Q�a�B�7J"���U��m��}��'J�'��'�^�@E*�Gx��G��(�`�*\�ў'���+�'���'�R��$(y>�Г��
���@��L�.[�=��>9���?QJ>1��?q�I��?�G��-�H��.�( ��({���
⮔͓�?����?�֑��ΰ~���/�f=`s��>Q���ץ�!�ԫs�i2�|B�'�N�#�y"�>��ˁ(�����Y-	��a�X��7��O����vT�d�On�O1b�'C����G ��_-n]|x�㢒��(O����O��;�+�O�O���1f$d� �J�?i$����^�6m_;S���OV0n�ן���ş0�ɴ��dٴU�H�A�_-M��t.�}|���'�⣖�H���|�Y>D�eӔ��"kҜ�R� ���p��i_B�aӪ�d�O����O�8�>�"kG�m���B��P� �@y��G>;��G�x�R�|�]>�c��u���I$|���W�J��ջuE�<=ݨ���4�?����?��8�'�2�'��*X{�ȱW'��~�"�Y�@�g̱O@��:O���8O��$�O��$�KhT���oV(�a�ʁS`�n�˟P�ɴ�ē�?�����2�>?���qjfr���u�g}R��U�r(��y��'�B�'y�'\�Ra&\%X3���1h�0et�QnZ��'��|��'��H(H����c
��|���"I�H�J,Cw�'^NA�',��'�����d>�Hug�#��h�gC#%�8��>1���?�I>9��?�Adڝ�?�3��quJU�G�B����@����q�����?Y��?頕��N�~��quTtcD�	�>ђ���h3���1�i�|��'�"%[0A�2�>qŭB2E ܨ�0#E�x5����)�Ϧa�Iԟ\��@y�X�I?����O����O
$k���@PAmJ*,����dDJ}�'R��'-T��S>������`%z`��*�-�XP t̕��Ms�C��<���[��&�'���'�0?)��Yj{��$!�I���(�Ȧ9�	ٟ��q�%� �O���!ܴYeX$+�/�����99�MlZƟ$�ش�?!���?���p����!LRxp�PΊ-Tԩ��iY ��?I��O��)R�'l����6*�p��odx�C�\�7��O����O����s�i>��O�uY� ڭ4���!o��[��5X��i��O���ƼH�D�O�D�O�18��L++O�ٛ�;Os�4������쟨�'zh��?�O>9�Jϝ+䵩�CԂ4�ŢS6j��'�Е1�e��y��'���'��s�����=�ّ�%G�g��m���ē�?I���?!*Otʓi�����N�)n��D��_�T��E�<a���<���?����,�j�S-�(!�/ƴ�p��itOB7m�<������?�,O`yQ��i�� G�]	�e$�X+v�<b&�������I��ħ8��ޟ� �,��j��4���
���9�MK����?A��1^���>i(W45��%BK��Iq$�尿�	៤H��v���	���	�O��$�O`y�ʛ�a�B��L�fπlQ�.k������)��#<��OS0���
G��Zl{�o��)�h�ܴ ��ϓ�?A�iz�'���'�� h4%AŦ`L�Il9H!ߴ�?Y�Q���Exʟnt�w�i̶����Z�n�9F�h�hD%NЦ��	��M����?���?�@�d�ebpD��xO��D�Srp�l�w[0"<A,��{;O��ė�&��li@��%3���Hl�������I���'&"�OX�M�T�mI�
5D`�}���$�?A�ߑK��$�OB�D�O���O�]m&�i3��GU���A�Qݦ������J�}"�'�ɧ5�	�$V��`����x�Xh �P���V/�~�Oޗ�y��'�b�'�'4�zZ���0��ܑD�ρW�oZ���'�b�|��'��-kɲU�v� (bn|�3��)Pɓ�'H��{�'��'�b���ou>	Z��V~*lpX ��	x�I����>A���?AK>I��?Q���e}hȐ1�؀uBY� ���'^~x��ݟx�Iȟ�ZwB��՟��ٟӈ�1���b��%����M�M;�����?1-O�,;בxR)�8
��Je���t]�4'b��M����?�bAT�<q��]s�Sן8����G	W|�1��E�|�D=2&n� �M+)O�ʓ5Bl���🛶�'tŸp��v~6L 6,�$�MsA��?I��?���?	���?A��?s��3~��hSa�{�H4��I/H0�f�'l�ɨ��"<ͧ7�v�o�L�D�c��I<BHE��j�F.V6M�O0���OL���OT�D�<�O�D}X���&.e��#㞒]fyzb�>Ѥ@[a����A-�y��'j����\�=�~��䜆k�*	���m���D�O����O
�%�$����T����E��>O��D#d�	#"A �E~�X��yB�'o2�'�~܂�o�%@�X�P*�.\���9E,o�����O�H&����ß8%��8� �uر�$X8��b
�3MN ��W����g�d���v���֟\��Y��@#.,@��ͅ@N�r�̽T��F�"�d�O���6�D�O��d����S�@2`+��3� �d�I ;O:��A=O����O0�d���ʧ�?��ϓ-"V|	��8,� ��tnБae���'���'��'��S���&Ӱa���ϧ
T�%a&�	?��������<Q���?��`�O$b꧅?����d*n�9�)
3�Y�l�=I���'4rV�ܔ'C���ɟ�	�����uɃ�[��mQ�%Ӂ5�Z6m�O����RU��d�O����O����O6�$1be�uA��
�쳤#�HA,-'��	ny�@��O�nZ6\Z��U�ܖ'������u˛fD���y��'�d6��O��d�O���NL~�Mؗ\�`U�v�_�p%�p�@L̮�M���?Ԭ�J�'��#z6m��S�����j�T��`śv�'��7�O����O��p�s�<=��"�hը�I�D�M��iż���D�|j���<��`.���s��!{��CP.*ohZ�i4"�'"�'�&O�d�O���:#C4�ٕ�(���H
V��b�$Slu��*ǉh���I埈��DV��)o�`l �A5L��M���?�5���OV�Ok�'4�5PB�P�j��H��D?&��� $&��	/��IԟP�	�X��.�� �+}bfP�'����Q�A�i�&���D�O�˓�?����?a��3�D���T�::���d)�V5ΓL��Γ�?����?9K~"F0���qE�1T*(�P�M�&{����i5�Iݟx�'4"�'t2a�.�y2�ʡzK2 `DjC(.��@�>p`�Q�'�B�'C��)��XC�D�'J2�	0S=Y�n򧞱nޖ(i��f�D�$�<����?��
����ܴP���Qh�#�,�%���ǿi�'�~C�'�Ҫ�~j���?���*��PH�/$eS�-�H�ZA�T�|��ڟD�I�]n��d�?9����%�}@��-l[ ܡ�f�F;O@������IڟP�	�@ �O���f1fűb�Q �~="3.�==���'W��]��yҗ|P>�"fӬ\X�HL{�\�`�\*�@Zr�i��oӠ��O��D�O���'���4p}���6FĶ, J�(��$ƈ�:ش<?�a�����雾�����g��)�ӫ���y�e���n��2�� �KbH`)1B�>Oܾ��R�������7�Sk���Rг�銫Q�ɠs���Y�Ƚó�
:e�����,pH:��4"O�p�wꍥM��)`򀄣Mژ[abA�L�(����yb��X���w8IR���;� i:f�M��$�y1�)#6������mJ�Dq� �!/�)�!���ХP�
S�d�Fy�%�L�	13~z�	D+^?v�T8rq�
w؁�F"��J�ʅ��Ȇ&S�УƯZw�gm��
��Y-&>dHC�۰,G����O|��<����?�OI�����N�jpC�l�+i��� ��Y�W@Ȓw,���k�� ���a����Tg�'�|ظd��* 4�#DM��}a{"e���?a�?(|̛�b�:F�� � ��e�8]P���)�|d2]#��&"������L V��ȓ����&��E�D	�J�A�����	cy��Ѽo"���?�,�Ьk3���V���ᖄ�$J�}[A<O����OX���#"�0j�F�`�O�]�f�`�N2*%���@>I)^�<fd[�j�&9*c*Dq�<	��L�
��4�@L�FVf02D�ɢB4H���O��?��aƦMe��K�J,lm��a�t��I��,)#�%WO��0�;M8��d≕X��1X'��3�0�萫F���?m�;�O��#���ON���O�P[����8Ǹ	�Uξ����/!����pN�J}*hJ�F��ʧ��?�b��7J�A�
}a ,F�&w�H�bMӪ~���p�Y+���񧈟2�05i���sl҂p I{��Js2S��'�"�����O"��#�y�Y�$��",�x�sA"O6|c���6��@�a��${��"���HO�өj����A�)%ƨ�Dˣ������)�o��M����?������O~�d��*������P)2lx�HbGL-P���ߎ�)`2�K����I�%��5P%[�H����N��E ���^������f��;ǓP���s �7��A��ڼi��T� sH �����G{^�$��N՘vN|�z����X�".D���B؃td� �N.P4쬡!J��HO�M��3��=�v���E͂��&��ͅ��d���Z���NX $��R�$���jYw$\
t�N�2h�̆�@Yb4[ɓ6�1����k^h�ȓ*2���w$F�a��I&@�����d�-ӕ�=xF�y(;H��ȓ(s��c���R%Jc�� ����Z��E�P�MX�"5�9#]�0��MWB�2Q�3��e�v�C�1�Ll�ȓ$#�u)E�+%i.\q0)�PZ�!��S�? �}�ǂ�z�@��B�	G�<��"OH����H���J$��3\��"O0�+�ăL�\�QT`�:@S��"O���U%=9�0D�6�DWU0U��"Oȡ�/O�XQ6��3E�$�H��"O0!Rc
��^�sD�8$y���"O�kw���m�L �C��k���2"O4���m�+#�l����{\0Q�"O�`�f0)a
�"r'�.kTy��"O�T�R-_4B&M2Q$�Ksʡ�#"O0� �I\�q�y��M	Ok��I�"O�|�E!�n?z���(�#j`��"Ot��	N��XQY-x�"O,����=k|@q�G&�	����"OA�$��6D؀��0��T��bQ"O�ؚ���bߜ=+�b^�8J��v"O�Q�fl�4�HY�uk�s;���P"O�u�Ba�G�� �$�1-F[�"O�5��	�&UR��D�̍ˡ"O���ˊ3	'T�	'"D:V�-�"O~��H�N���C�ܫ< p�1"Ozr��/Xx�}�w쒒&(��y�"O���ǥf��{��"��0�"OHi���̗�.d���k�F|C�"O�e�&G	 =|�;����k��5�&"OT��V�Z�yH��2Ԧ�r����"Ovx1bN�wHfI�#d�o�||ؔ"O���c_�X��ɒ"I��
<�C"O`ii�f�F���e��"��,�2"O���B�6�����I0h��yP�"O�}���r�����݈c���#�"Oj����=e�(�0gҭ=�$��7"O:���o� �S�X��PU"O����۲AcT�q��g��!"O���E���o(eᔣ�mnp���"O�I1D�;a����́1<��Q�"O,�[�fό/��'+m��yA�"Op���i<x��Ui�j������
O�Y��CV�n�>�ce)�W�t%�W�2t��#�^$�M�%)�.���k�`����	6����{�H[�N9�8!�!S�W�ye��4�yRAZ�.���F�8Î�ꃆ����It0�=ɍ}��@J�z���(�j� L�.�y�@)��(ꔡ��T����Ыی��'O�T�Um'O Y�G۫9	���Ǌ] (M�
O����<=B5�j��N	A��7>�\���}Ȕ���W98�H,�*�[qN��	Z��(b�{�ύ,:</���1��ȞX��EX�'GV���� �lUQp#L�8�Ν�N���"�G��ا�O���2�nU7#���lߍ-�	)�'8J�a5�A�k�.����L�}��{҄�"����dP<F�H�d��Gm��0��&O̡�$�g�ТL��4����\� ��U� o(<�剤����F�=|�l҅�Lj8���#���'�>�'a�-q�V�'�H�5A�5��'�v��6HO�_�Xs�Β(1<�XL���f���اu�{�
hM�p
�-Ҫ�R�L���yn�:Y�*uH�EH>��X�+T-��'�x">+U/�y"���Āh$��<�^��)N9��xB� �h���@�d_�6XJ�5S# �\�=1+[=��O�!�%�ߙ=����P��!&1�hc"Ovu�/��(x-(4(�b�h��'���� �'���G�D�xƘ�7�Y%=T|P�u[�u�O�� �-1��i8�m�O"(1�"O� X�F�f3L�YfL�z����C0����$�T�d�W�9�`�k&b��n]!��3-��,�g*��$�tH�!�7-����)��<S��K����S��J4��F�`�<���ʉd�����O��;�(�_�<�ꓛh(p "5� �Rl��MR�<AE��9-��(%k�$N6�rqO�<�!�*�Ԍ0p̉�u&�&�Ay���3#�a|�"\�Ws��[R�En͞��D���>�vD��yb �a�q���ZY�8󒦙�y�%�Mo�U�T�b�R�����hO�Q�&D2�'�@ ��[j�d�1K�S�XĆ�[�U���m��9��
-^�I,2 ��?E�T�A�h�����o���l��I,!��/A�(mIp��HZ�\��K��;�ɇ20I��I�����ČK�2X��ѓd�>B�=F�>�Yr�֛��rJ�K B䉐"��!w/������%�mp�C�o��%��J�"�^t�R�M�P��C�	�wi
�J
�|*|`��̯
��C�I�[��8ԤXT\$Q"(�u�C�2u��t��׬s}R��D��%D�B�I("�F�x�
,8Z�I��F5k$�B�I��
�8E$��*L�ir��'g��B�I��Q��/�/3xDa"�e�y��C�	m���w(A�A��("�X�!M�C�l7]!P R(\z�x��C�	6E�@Sq�Q�v�p�ӫe�*C�	tcMt�:nކ0��	S��B�I4��w�ʝe1��4��`��B�Ɍ|�4��Hx��	�!	Χd�B�I	Ht9C�χ�nP*A{�j��BB��/L�6U�#��<�V|�t�HhTC�	oPx	zE ��):�m�e#��8C�I,�F�r�m@�������X5C�I�3]|Ax�	P$$Ш�Z@�պC�ɱx�t]S�*��
C�yC����.+�B�	o;v���ٰ.s,`v�Ѩ7��B䉀/`���,V�h���`�(��^�|��������3Ѫ�(�M�ȓ91�mˣ另G��Q�S�/ 8]�����X�
�> �ܨBJ�6|f�4�ȓh�����o��r��s(�4o���ȓV�(u��׻f���j%߸Cј1E}�S%=Yj�+��]���Xs�QY�D�	5�F�"BNX/2HQ%��b�NY-6Xc��>�8R��E2lrT"� 
���E���`�����@��<?E��K��*�J�m�Pf��7j΢�Y�I>Y�jϠ�����!o
Rf���o25r���O��]�'�:D*d�.A�U���O� R��!]�4���őjIJ��$�x8�H2\O��Þwt����_�"��B�K�Ƅ���N<8<�u��f�7M�#e<���O̩�&��W�~Ũ�AA D�ؘ�5�ɞnc��;��V�^��F���K9
K`�SЫ
�3"٘�����'�G&o�d�!0��FW�S�~2hT��F�3�J���8���I'<B�	��E$"h��S�84v4���G-_e�,����u��0	[�6������؀(�� e�m�ܳ��O�Ÿ�@�-���i�$�� ��	�jMr� $Ć��5{z����' &*��#c�5PL�(r�Bc��q�Ә?:vxC���Y1 ��>��M��X/R=\<nZ��QğI��A�O�IVT�6h"Ο�hQ_:����G�����o��y�L�?"9�N�?�D��7G�c�̕�'��`P��7D�:�`��["M���)��f m "�ҲmيqC��D�	��z�dK�"\!(Ui��xZJ��r
M L\�q�c0kҠl+�̀j�qO����fAw�g�$�g�m��_�_�4M
p�B�&�qO&�R)V3?ٴ9�f˘�c?���5vU��)�F�y��
�˝<n��}#��hc �+Y?ML$�$' *,�x��2�!A;�����T�	��l��H��)� "M��lZ������k�=49�q"f"O<�"�K��Zx����A�9��`� �i�z��R�r�>�8�4L����M�ch��X��\�u�J�g��?y��{��;֜��C�]�#���A����}�Z蔎�,%�p���<�Px�h�_|����G,>;��������9E@L�烟#z���?���k޵[�h �F,)� �˱�7D�d c�Ր�,<��a��̭�'��OZk���3>��i&�"~�[���	!���0e��y��KD"O>�p�+Q��Y�QҨ�U"Or,��� � ���Z�6Ȥ��""O�x3%ƛ*$Q~�kf�ũN�� �d"O�|�M�6[p�	�*�k�l9�`"O�i Վվ2,�m	�e���ö"O\!S��(tX�A�An�l�G"O�y0�͐�v�\|wT>\�!"Ofx(�b��;��9�oZ$*щ�"O���,X#I� �r6NѣF�P�U"O�X�a{������O�& ;r"O����׭.
4B�iF�L�d<9�"OF�b�nz�Rɸ��Pw�|Ȃ"OVa�FI�o����׎��@���f"O ��T��$'V��:r�/d1,�"OZY�Ѥ@�_Z¬×�!&��i�"O���� -p\Z��TQ,Q�R ��"O�0�e�G�&�4��A�!]t���`"O���R��ʲ�H�!˷H?�\��"O����>AHdȔ���&�=1�"O3���M˲�(�Fԫ�h)��"Ot�����ۮpSD ��Zþ@x2"O�Y���J�t��!p�DS�AS��hF"O*���!$���aUCJ�f�Ni�"O�da���@�L�03��4�f@�s"OVA��
E������Jl�Ԩ "O��t�� I��W��	?�v��a"O�d�d&�s�T  3�~��"O�p��ױ�� ɦ�_�g$��+s"O�`�VΌ�1�^5�BD�5f@��"OL�`wM��^�HK��Yi��q�"O�a�!�&����+�R��3�"O\�ڒ��8)-�"�'���c�"OXYA��[���LOD1x���k�"O�u�q�� �E��M!g�\X"O4]HfiA�^궵!5��"3v ��"O�5A�ΩK$�p���\�x��"O���+�lS����t��"Ob����&*�ެz*�.W1ʳ"O�T 5�q 5�H�s�Za�w"O�`�u�
%yἼx�GO�YB���"O��{�JR :�ȝHtF�+�\� "Oh�a�C��U(pFY�<z��"O��x��	�>�P*1�Fm<<��"O��S�Jd6%�U�OqN6m��"Oz��b�
L��p͎
3B��6"O���F�,�|���̅��؛�"O������Pt���we�8p�� �"O|��H�{���6���g��z�"OjIN.S�l���` D��6"O0(�D�P��]����@��I�"Or4�4��'2i��O���"O�P��ޅ/��%z0`��N���"O��
��L�Τz���)^0(�"O� ���{���˷hǳ	ԂT��"OBY+��7��5��F¡63Pܠ�"Ot,�c�!jTJ,㥝���q��"O� �|B4�ǄE�ؘ2eJ�G���"O:��v
R�
tmC�4$�B�`�"O<4Q&F�U��Q�gN.Iz1"O�MaW��c:����+��Q��"O`�IPJ#|e$@�0��LS!"O UK���2n��[rK�� ���Z�"O���#���:�6�*�7 �#0"O^���L΃} cq#��B�� �"O��!eI��;g@��#K���[�"O���A�ܠ\����ADh��P�"O�8k �J�|���rւZ����ia"O�Թ&	�.�V��T�B�+U"O֡p����AR� �#$$��"OhD)�"�3����b@��Y�̼!�"O�p��e��.>�0h��';쮹�"O�ԁq��u���m�q�^A $�'D����Jٰd�����6ihn&D�$;���&e�)�G��*3�Ν[��/D�|�V�Z�zQ��Ӧ
~�iY':D��!2�Z2d��W&E�A=`��<D�8[ ׀F<�d�W�a>�AB6D�dґ�I����7�AR* 	�S�9D�h�F�W�~0�F�I6��SW#D��)�D��(�h�m�Pj���#D��4Hլ<�l��A��|22B4T�$ �
��(KoC����"OrU��ݦt%����"\��\x�"Op��1J��'z���Ơ_�R��"OV좤�	���AR�v�YC"O�U���)�����?C�hL[�"Orx d�"�q�]�L�葙�"O(x���F?jl����
=%̚u��"Ot(X
�	1��H� D�`"�yK'"O�IӃ[3<��M�`�P%^A�z'"OT�*Ā�:[�����>���"O~�SCL4R�� �����!��&"O��"��7^��d`���e�dܺ"OְZ�FЦ���@�Z��b"O�ᐅX�`�с6��_����p"O*�R/ʳ#}\$J���&�05"OlT��b:p���!��A�/����"O>�s��ƃE��9btA&3o�U@�"O��R')�Ƽ��Ù2K~�bS"O��;���c*f����D/c6�+u"OZ�d���]�`�9dInP
R"O�4�DµX��p%X>u3�P��"OF,��`�@�P1&���<*l���"Oqs f�F�l@�c逵&9�#"O¼s`*F)ch ���- �"%"O*p��J��I�f�2^��a�����		{�4�UJ_����J��{I\B�	�n&8� T4�8b�^#;�C��):�4����! q�����DFvB�I����Ũ�?�v����ƶA��B��k0��B&�A%+�t��a��3�B�ɦZŰ� fJT.SDu��,se�B�I6bc����G��aB5�ċi*B�	+kf5BR O��˓f�44�*B䉣Q=tmXe��|�aZg���C�I�f��Tȑ���gyrA�v�	�v��B�	�Dh�<�7m��i7Jq��IS�rT�B�I2�~�yԙY)��eO46ϞB�	-I�6����@
&B���{QtB�	�j6�6'F(6����oS!`�NB�)� �%z�I�{�M[��]���B�"OxI����LӀ �7�7�*K�"O� RcU�zeZ(qf�1��R�"Oz��d��-P5@�$J�>9��"O:�ãO٤M����V�Q4o�t�i�"ObPrfcx��'$�y����"OB��vO��N=:��e/�a�"Oz�A')
h�Yb`A��)�@�"Ox%��mթ^(�rG�x�Y�"O�,��)J۸�Jd�^�2���r"Of��ŤWc�i91�Q-y��u"OJ8�0!	`e6�Y���!c���G"O��Za�I�	 R�J� ��e+�0I�"O,���f�
 �̅Q ؈w���:�"O,��N�����k̖�6,���yr!�(}�� ��U�5,l��&A��y�DL;=���j��KVU�4pw!�'6]���3BB�����,��܊�'xDP3����P����.�+���ʓق5���S2	�h��G�<c���ȓBn��銉5�:h"iR�3�^���m������(fp�1DM21��E��l�B<�MM;36q02�O,Vh����.[�*WR%~���PȨ=n���ȓ�H��� �|���qFg���XՇȓ��x2�i����ă6]n@�ȓ}��a��'I�Z�Y��ɳ�4Y��#�&8�&�4��퓒��J����=�	�.������J_$t�q��0z����ȓ��H�B@�~���y�/ƪ	�Іȓ��D b]��	��������ȓ�"�*U�_9"u��FI�5�d��ȓ �8s�+��[�}��'�|+Vن�Wx��1�N�nT ��@-���@���F�p�!�����N)H�<��ȓR�J�UoD0T(��R#)>n��'_`�p�"AtF�"V����Շȓ_�D��A�#:��d�`i�4����>�����T�xH�eMΛN����JO/�y���9Nr��sl�@z�T�f��yb��*-9%�,H���僬�y�a׿j_�أ�j�
Q���X����y�%Hrd-P� 
]}l�2���y���b�i�GHI�UҠ��G�J��yrE�8e$� �RQYҴ��y�K�;1Ԁ)Ս7��lq1�Ě�y�� \j��r	�v#��f���y"-��q�X���͔#,4� �
Y��y�ޗ[�VA�BE�(�j��A@��yW�b�FV.��#t\��	� �y�J��x��ä�8Lݪи�M���y���~�Bt��Q��h��G��y"�
�K�LU!If�	�)�9�yA�1T<��ɉHgv%�#M�"�y�揣6��t��<�;�bX�yY=({�	8���^�T���F��y� �qN\Ѓ��W�� �����yr���x)�m0��"F����DaC	�y���zN�u�ӋχC��j�gW��y�d�<z���q��X#;1�3�Ó�y�Jic �X3FW�^�	�+�.>��|��	6W��ug	��Mq�E�NQ�s��C�I�$��p��#ǜ����ԾXpC��p6Q��Ԁdj�uN�C�C�)� �ղW�D�L	~�p�(׋Fm��:�"O����"[�:��p�d�}S�q�4"O�ub��/#�A��oX�g��tR5"O�qaB��r�2�B2H��e���2R"Ou3�↥�ݺ�g@�z���"O��Pc��j����%.Y�B!��"OZ����Øn,I��"ƫ%��͑#"O P!cN��Ry2A���J�l��U"O�I��
8 	Ԁp�-��1H�"OA�� %��-T�/0h3�"O�L�4s����鉱@�`�#�Q�<�q�׼T�n�k)Ϫ���t"؄ȓ3�~I����$r�X#��>R셄�v�%r�ϔu)��އEm����&\��V�$y�(��Y��ԇ�ͥKz�ʔ ,��d��U�=D�@0V�J�TnN�B�]�]��=D� 5��1�e܆�K�j:D��ɣ��3(��a�A�b��x�'H�R��{"�y���;Z"^���'�(J�h.g�VL�N��:�� �'|�y�'�:JI d�D�[�$��'(���#e�w��La�*�gRN�	�'&8�Δ���-�[!Z���C{�<����!�����*��a�@P�<9�hE*;F���2�
l�XA&�UN�<1���$`�4�xC���%�nt'�K�<Q�"]<cv`�����J�V��% I�<���-��8��É$��dab m�<��Ɣ;'2���/D?p��e��f�<QC+�yH�#W옪�te�%
�a�<���(V6�#M
�uX�d���i�<Q��R��-�Z
�T�N�::�C�;s5�1��e�	
�a`Y�C䉃G��ypc�x_���b�����C�I� ��+v	)�X8k#T�|�zC�w���N�Nd9(q��e�<C�%�2L�dY�5��܀R$D=\�lC�I�'���N�q�X�)hB�\9�C�	�v��PD�kՆ�� l�:C�I�fq�ɳ�%�9C�Z��*��<�XB䉷>����E�@��@6l[f�C�#V,���)V�T��	��`M?3�B�3G �@�S$Ə-���s�4c6ZB䉔'j(��0J-[���a!?y8B��^��zff%�ܙKB���B�I�Y
��u�	 �~��M <~�B�I�'�}�ծ�e��`��k+U��B�	������I�| B����B�IB��DJ�J�-8�`%ҹ<'�B�	g�|��a	ǘ9�쩺tot�6B�Ʌ/Q(�Ȗ��82�ٸ׎�>2B�	#H�(!` I��T��rb��l"B䉌%��3��'%<��$@9DK�C�IN熩Y4b�d2@`ؖMtC�I!8�u� jd�K!��OI�C�9X�E!֡�'0x��nM;4(�C�	���\KU�&yGB��c�2N�C�Ɋ������eP�+�,��hz�C�	�RO䑑��i���!s
QKDC�I�D �!�����1(Ә>�(C�I
P\�ħH�a�o�4C�ɾ}�}f�˓H��ÑL'm#�B�	A�(��q�%u��Xd��y:�B�)� �ѱ䎊>s�F�R�N�I&R�9�"Oة��;?`ب۵�](���"Oxuo�LW�c��?7�u�"O�H`B �/TP��B�D��U��)"O�$��TJ�fI_%N�(!4"O,H���xٰ1� #�Q�"On��'i�2K�� �A�Ew�T26"OeEȃ�J�j�����b
���"O6��H��*� 1�!�0D��s"O�M��M^
 �eZaGY8Q�i&"Ot��f L�K��b@�Z�j�fX"�"O�m�W,��82np�F��K�Zi��"O 4 ঐ0ܲ1�&_��F���"O�b�z���ӥk̈���"Oz1h�&��K�.eqUkͮ$,h��"OE3��$):�$H��^�q�(d��"O�t����
O"9�tP9\��Tj2"O$��6��<w���J�MUsJ�["ON�j�园BPj�*6"�l3l���"ONX��/�.l���!�GG(&���"O�YSiΠZ����ƒaFn��"O�M��H�&?@(��˴�0I`�"O��w���P ���r��7"O�!j�i�~|ʼ!��ޣF}41�"O������$j�XAŔ�bF�y��"O��A���&���B�ʰ1�A�	�'���Fȷ;d����ℓ�L0�'�d�8SK�,lfH9�)Y�w�┠�'mz�AA)=QEM� �Ϯg��Q��'�L	`�C�U�\05�Z.����'nD@�vW;�����Y͆���'�ĄQ$�Y){�H����T/.���'
�0
r��MIT�ˡR$�yb�}h�p�&C%:W������/�yMW�.y��+82̠8!(K��y���SX�ဎ�'<�X0o^:�yr(�"J�H���(�	�5#�l_3�y�×4�(�Ԭ?~ԜT#C��y��F�(�4	Z�(�q��(�7���y"hE�y��xCb��=f�,m����(�y�j0V
r�z�iҚahH��燅��y"$\xW40�2)�<B�䁘G���y��	�0�2`*�
�h�C�C2�y�`;�69�7&�j�Z�rS���y��O7�b�Y���+`���Sd���y��ULYsw(U?_W�Ԩ��y��?Zq0
 ^�|u
!bW��y"H���5;�GCv�e��!�y�	�iOv�p�
A+O��C%G�y��R�\�v09]ن�q���x�6B�Ɏ_���+�A�-HJ���U��6h�C��+��xw-�%ab�򉈇=C�ɾO�L��L��_BnD�5)�\\@B�I�K}�|S1�N]{T@�ؿ"dC�	�-�M0��\46�,���F�RIDC�I$GON����0fRݛr��C�	�f#����M������é@�C�I�m�ԡ�f�05���Id)�V�C�I"m���RL�:<<��%*�B�ɩm��q�i);� HEȃ��RC䉹%�N��.C=w�X3�.�?U^�B��4S����>D���Jc��B�	�$@��j$�ާ
غy��$��cRjB�Ic=\pv!��l�rT�@�JB�)� ~Q�+W�k�ypc�1rd��@V"O~��/)-2Tcd�B�Z9���4"O �a��^���rB��!M���5"O��2�
�F�B�5/6���"OH=�G	�v䨜���ɯ[\��"O� �"X�	���R��
= ��v"O,LK�j�-��%PT���:��t"O�0HA�&(����?ZH"�"O0$3��	�N���qe��k�`�2"OH����%�ŋW�M�Fl���F"O,��eY���Nόq^���"On�cA�,t6p$*���f7�ظ"O�|����'_�> �Qq��HA"O�@ �F���TI,"�B���"O��R�d��SL��Ӥ� ��pP��"OLT�u�K�,��!q%��=F�
��W"O$X�!A�DKfqcԃ�1g���"OƝ���̯+}��PVBe�$8R�"O$�;V/X�(TNyR��hDA#"O|l�d/_�4zi�d�َ'�M��"O�4��Nޱ<p�1��<_�PŁS"O�!pҢ$�|٠'�\�_g���"O��!�'�{6��2a�L����"OB�8E �n�9�T N7Q�8�"O��ZRȟ&	�`8@�ϻ	º��"O�̀��F i��W��%̲�p�_m�<i��	��P��@Îp��e�Sg�<Q3�Q��NDz�"�^=$���@b�<�3��O�,U�,˂Xd��u�b�<��+�91�A�5��v7j�Y�H�]�<�d�_
@�b��`EZ�x�|,�� S�<�ÏM�!��gËc2:��$�	M�<A�o�	:����ÆI��z6KK�<�à� %�!c�� ~�&*��I�<Y��ߔ("��!�zf<��6��m�<�W�m8���3d A��l�<11 (�x�+ՠZ�\7�5��XA�<Y��#L �Y�aM0	��h#E
�|�<��޿vp�p��/�Jl����@�<����bd����R�V4u�z�<��Ȋ1�40�m�WRl�E�{�<��!�7N��kae�B�P��D�m�< f�4k����NB�*��+�s�<�����������Q�/�r�<�"^�z��� 	F5p��Avo�k�<�@��yW`�[���3(�ڱ�m�e�<��%@[��0��.�t��p���\^�<�uf[�V�PL��nN�Ce�kS^�<	�B�\� dK�1���'��[�<�V�̞T���Pm�"�h��pd�P�<��G'���8�J��v�
e�"Se�<�s��l<h���̣{XH��#�w�<aB@˂|w> y��� w3<�⁯Em�<�g�вFм�p'D rc:���I�p�<�Ϙ<*��"'k�0<��12a�Vj�<����>�R�C�FX�t���jIj�<�iΉZ`6�c֧N$8�)tL�<e�+c�f��4"�R���*�l�<�rlH�G�zt/�9S�	���i�<q�A��C����,����p�Rb�<��g��/���h���,�x��5B\�<y����d~rx����6{��D	Э�~�<����;G¶�!P�Tڪ���&�w�<!�&�LȠC��.p���g�_�<� rT dM� *��1Z������"O����N�p�,8w
�s�v���"O"hx����BsDqj檅�lr$��"O.99E�Q�"�`&j�~n�U"OlL���������׬F�)Pb�F�<A%�S99@�3�3� �9EDA�<��*"-^��`��rԻE�VD�<1�NF�[�������2�~@	�I�<�Ҝdf���L� �|�[�o�<Y�!����8 F��y;6���O�<qB�(��K��E�L�PX�kr�<I�e�"zSJ��N�w�8qQGPw�<	��E6&|��2%��H>R�����u�<9���m� y���F�a�+�v�<!��}@<P� �<B~pq��ퟰD{��	�%�z�q�-�h���0R�ߚ&�VC�Ir0�z5f΅N���x%)+I�JC�ɂ,� mB�U'L$V��&�t>C��R^���5�RI��N�~C�ɼs�D�bG�h?���)��B�I�H.�d�m�*.�:P���W� _�B�	�|	�����lKV�R�S�0�΢=���hO��A&�J�� I���y,A#i�O��tG��'9�5�U�T�\pS�Nd,<!��'��p�F��_�D�Is`�`m��:�'�H�!$*Y0Lk�躒"ˉbF���'E��C��g��uz���M���	�'�t��F�߿�$M�Ej]�Fz)��'��,s��ޮ{M����lC)<�z}!.O��=E��܎]Z�(f꒓<�@��,K6�y�(o�Y�G�O#��l�QE��y�^�{+v�q��N�0� GR�y��+�������dM"����yr��%P0;�+���M�?����Ӓm ������!�����2T���c�V���Þ9}$����̏'f�`&�0D{����(oZ"7���vĨ�$���y��e�4i�l�1P� �@ �yG�X��}���l����Ǡ���y�GR0 ��t�5���1�(���M�+�yrF>Dl��#�,T�'�A���,�S�O���k�I*g����0	�F���J�-���%�����s��!�ȓp���N��Z�s7�S��U��< �12�E�-��e��h��g1ؙ�ȓ6`�#�!�x=yd	S8 ��8���ҥG��hɚ�FmM1F(���ȓ��ES�
��D_2-S�1EU�P$�tE{�O���'�F,�d�+v�ا�ִ+BB�I Th����E�J�zx3������d+���3�V�l2<�����soF�s�e.D�l1e@�8��b@�3370�,D�89�	���tqx�-ˤ6� %�m'D�4���P��@1'H��,����7D�x�!l߼^�^ ���I����g4�D%��?Q�ON��v
J\z�-��
ع��	�"O�-i��2�^�&C��T9���F�'�!�N�7���`J�
X0��+U͋b!��ņl�Lj#H}���1��Z!K!��j z�A��Z+�,m��j��4`!�P�
јL�UF�J�>4z�*��gG!��7�"$���$� x�E��@!�Dʜ,�� ���bpv�j��Ɣn@ў��,��uP�˜$rh-+�i�� ̈́B�)� ���㍔����ǌ._w� W"O��SFL^�`#����@C1~hY`B"Om��(��G� �@-���2"O^�����)����D��>&��<��"O*h�@�4|�r�@P��)g^*�"O�hx���9/�ѱNE�R��|�)���4$nҢ�@cN�c�W>�h�*O���dh��+"��360�(��D�Zc�%D���K�"`6PHU��
A�
�J�!>D����!f֬���-z �r*D��`&�צGe��ńL ���'`'D�e!E�����w�l�Q�%D�|�4�\1@5b�k�
���� Q�84�L���b�4P3&�P�.ei���wy��'K���&��Y)��I�A�a��-!�B�N��!r�<M*�c	"�B䉫DӐ��3�6i��#	�nC�I�m�B�#���c�n�D#%hC�	-�� ��$ �z�!�&�2�ZC�IjB�HI���1.�j�I�\���ȓd���0h[}�|%�����e�~��?	
ӓd��󗦞�U�Lpj55x��ȓu7~X(%`�j#�J)N֐�ȓUw��c�JQV�x,��g��"��	�ȓ9����:UJ��q�\�-~����L<�7�	��D��&+4�ȓ2Z�]ӤZ�qQ�ݙa��E{��'�`QzUA�OB&����%�|�(Op���٠#V�I0fb�I �ٲ���!��;I��pe��D�궬��V!�DϷq�Dy��ʉ)p��t��1#�!�D�  �"�E�*U�i�eF�[�!���Id�!i��1v��m2q�/���Ο��?!���j۰�j��a�8�3gǁ	�?I-O~�O?USe@_V���[�,۬TʔP�taf�<�H�?מe�h�&s:,+S���&��F{J?��NSr�T�:b�s�F��k4D�d#�^�?���H�葾n��H�q�>D�� R.9{W��f�a���@ <D�P��+߈� ��@�C^(t�O�<��B�0�� 
d�0&���S,p�⟄�	L���芷j�PݡS�M�.��]���0D�d���Ѵ|�pLi�ʴRK0)+⬲<�+O���d�,d����T�\�C1v�J��_,<0!�AH�t�22a�9]1��ɶ�Q�7�!򤋹���A!c��o;��ar�Q��!��Y4w�|T��΂9-���0��)?=!��¾Tɶ��'B�!�u)��ǅ4!򤝶3��=����Y�
�㭐>"!��B7ah24�%��3�Hl����]r!���"e�*qL������Q�!��� hk�pY��f޼����Ģ`!��c-��`5��5r���x@ X�	!��W:4*9:�gެI����!�$\J�ʠ�bIsp��P��؉m���)�g_XZf���Z�K�ɉ<�͋�'Q���%bO�Q�����$�&�v���'xP:��Թ!��@6�:"~�9
�':"Yy�,�p�dMSuA���k	�'Q��g&AT���#�B�W�d��'�l�H�L�.g�ֱ3�f�;}l-"�'��ѵG�-�
��$w�)
�'�\��'픞B����7ț)t���'G���*� b�Fpa��F��L����� ���2
�@ǭf�$| �"OVԀr���:��<:6��"O2<Ȓ�.��*��W:c7ؤ@�"O�,1�aI<< j5��7� 5��%�S��M�6�4��@L�/}��4�v�K b��'{ў�>��Ƕu0��׀�a�ܽZƹ<����	WC�,�#B�*m��`č	�xZn�ȓh�Ԍi��@�B��R��4br��ȓ/�|hs�ƳA"XhFş1l|:=�ȓ��r��%*�(�gői���<ZȊVĀ�a�V�S���
�%�DG{����B�x�02GE�(sXHy����yb,7\��$����pV��B̗	��<�����	X|A��t`���&�Z<6�'6a|�(�� �~8x�l�3<�@�F��y�F�)!� �0�Ɇ�;��I�\��y�.�]�V@a���6G��S��Ƒ��O�#~:$l�,/���Rp��[Pu!��	m�	Y���O���'c�6I=�Jr���+R�l)�'e�P;��I���9��o��Afȓ��d�O0�4+A��>>f�����v�Qx�Ȃ|�IN�Hr��D�dU�&�A�^�	��=D�Dc�K3Y\T	!+�	O7LM�3C'D�䛁ψ� ,�I�3K�<���&����l���M����i���.�|�r"O4t�bƁ`c���-�#n�(rO��6�.���R��`ExQ�Ox�=щ�IY�FP�����F�cD�fv!�$��E�9�`�s��m�F�3_!��S#�4��/�J�ci�#\s!򄚊����� �I�t�Zchü"^!�D�pO���"KR7)�؉KW�V��!���T!��n�w��y�C�P�!�$�*8(� ��AQ�h��$��"2���f�'�ȭ��G�:-<�`F��e&� ���'�<Ћ�d��\��I6cbY��'�P�T��DZ:�`A�*T �'G<���D^�v�����?Qdy#�'�D0��I�`�D\Ȕ�F�3Q�4����hO?A�R,���Mj��' �@DyuY�<A0��%ZטY)U�U�Tצ�Ŭ\�<��Ǒ�����)|9���p�	e��"��
YЬ��%�R�yE�6D��8P��8��� NG#8����0D�LHfd��y�TS�G	k��X�&`<D�l��J��D��"r��z̄����9D��KD��;@}�X��d�r��`;D��t�^�Fi���6|��.D�+�+��l�̲� ˊXbM��B8D�XS�[Dz&�j#�O[N��ҭ;D�к7��&$��\���I<l0;D�ȃ�#D�=����,wjL�`&�7D��+"T.t���!x0`X�`:D�<�b��"��-y�Μ�'����g�9D��P��*�Z%�M�r�x�H�`9D�L�6�	 l�8�gBF��`��Q*Ox����Z�J��e!�r�P"OJ���`���-�ح��N
�"!�®����ȯ,�@���΍�`!�W;�,���`_� ȸ@q��Ӕ3�!�Dǻq���f�����$��X�!�D�^��|�d'�%-:�|3�a�M�!��0*���H�7"@f�˅GW!���',�I	� 5uR� �Ìڷ B!�� 8\��\@�Qq��I<D��!�*O�%#G�]&@-N�qՇC�C��U:	�'����� Fd�ճ7N��U*O������7�*3曨
� i�2K[�B!�d��]AX(z%���F�,�� �!�dČs�Г1��!|��[�	�E�!�dM�8��	Ёì+�@(�5FA�@�!�D /C��5Q����o�j�3�
3c=!��'-��hV�Ǻ�D��.3X!򤑛�~ �����X�>�z�,�0�!�S q�9�u�ߩi�zx��(Y�!���֠�a�h]�#���`K
E!��9D&1XF�����jA% �	�O���$ثu�hr�-*�*����~!򤅊VAT]sfg
�b���Ǝ�
!�$�� r��@#�M�@(�df� ~��'�ў�>u���v���H��u�vh�=D��+�Z"�\�3n��k\R����:D��Pd��	T�ЅӆHN�Z�x'�:D�0������I0�9�"�fH ړ�0<-�2j���P׶ �A�L FB�I�P�=�2��r�{�ύ1f C�ɵZ&hsQ@	'눥�ӂ9P���F{J?� 2�'8�Ұ���X���d1�� D�<��I�kM의1.Q+92�ܨ�j;D���LD��,1��έh�hU��e;��0|�T` /d���S�Z)�$:��]�<�2�N;J�����H��~̙Kn�m�<ღY2Q�������H7���"_�<i��������)"��z0m�Wy��'��OQ>)"���V�@#�ƭb14M+q�&D�\��O� /���Swl���aª/D���T�W>���z$䓧~����w) �	Y����>���Ua�I�f!��b�4$�˓�0?i�iS�ctz����©�����o�<��Ú
F3$p(G�pE`�����V�<Q���G+B��ĭ� d[4bEg�<!P��1Jb����I�e��M���b�<���>�0��V*ѨF�����\�<�gO��o̖�)��_f����JX[�<��i �%@$$YVGQ+S�R���k�	H�H15IB!v,��`��4'�M�D!5D��{E*��x��%���1�4o74�p�Zy�<36&F�l����V�!���(JQ)�G ~slq ��TJ�!���|^6�x�ɏwZ�m��ˊ�F�!�D� N�qA���K��X�7k��=�!���c�Ԁ��X�P����IV
�!�D��x�8,i�PB
̀k�'>8L:�Y�.# U�6��5�ބ�'����"����0`���}9^	�'��{�p�"��~�"�cU��+>�>Lє�.D�8Bd�_<Uh� ˍ`�b�X��.D�,3rfX=	�:��!͝4:�F��&b1����?�&��Ș��8:��&dn����_�'D Pq�ݽ	uZ����5gD�;�'��T�%�ژB@���hʢ~�V�"
�'2b����T����G�]�?6h���'�
8�aЃ%��(K�6�l!y�'��:7�ևԨ�;�b�4��8�'JX��Fπ�2���ꀼ��@���$?Oz�����.��$	=V�`�R�'��HJ�"w�8�Òo��#�`���/>D��HG��;7�z'%1G�p��6D�� �0EO�hހZ�`�5�}P��|��$�O�b���Ҍ'+ܜ�QL�,"48U�0D��8�)�-�R��j�:Nԅ��/D����Ї^��pm��XL��.D�<�S
F�~�p]c�,� ;������&��0|�w��F�J]p��̂('nh14&^�<�Nڮ3��uU��Xc����KV�<)���t�J�Kg�?�����(SX��0=i��=^�5 �ߎ!�hd�7dp�<	P��I�f�[��G��-����p�<y�*�<!O⑨��� �����D�IA�S�O�R�3�	%uZI�UFU�� ���'&ў�D�D��`�t	�B #�.�S�"C3�y����5B�0CanP�*n� �ҷ�yR�� 4���%�?)��4���ľ��'�az"d�(D̣f�ٗL��@e"؂�y�e�Wa"�����v���b�y���~���ѲiX ~��q��M�%�y�K�aN����@�l�<E ���yrB�5���	����d6��@`F�y2�ω���j'W+(��wα�y�e��5Ҩ�J,�7�9k���'�azR��*c�Q�D�5Cʪ����.�yB`�V�|���O�#7 ,�VD^"�yr㘑]"@�v�ҍ=�֥��NS�y�ڿ=TU��&:��@&����'�az���~�SX;:A�,,�y���L�Դ�C�I�6(� �DD��y�&ϻ($�HB,H�2�8�(�� �䓩?�� � ����/&~��=F1����usT�h5eQKOh$QsA	=�\4�ȓ814i3)j�l���kَ��V��AD@�7Ը �4KԾX��ȓ%�.���^�+^���$j�9:t���ȓNT:A!1l��fl ��8T��ȓ �l;�b2Kb�7�T�p�jy�ȓ
2��Ya��dN�0��(J����38\!p��yFb�B���!Sx ��ya��ҕ�$�Ƒ
�α?\���	f~B��]ֲ�(f	�H�~5ۦ���yöun@�ÆϞA<��{�MN�y�`M
 g�UQ�38
������y2J@5�hB�l��<��K@��y��*r(!f�>I�a*�	O�y�˯K,�}8�-;=�ΝJB� �yrbZ�%�@ȕ��5�&�rB
8�y��I�J�� �c�(����H��yR���DL�0fƴM7�#����y�+�p;HU����>x�SC#�y��3ά��!�6)�$49A���hO��ĝ�	7^�y�G6��s6�Lq!�D�L�
	GhX#n �˥�� Gp!�$L ���'S2e�lȡXy��"OP��s��E ���ڲ`t���""Oh]�GC�;\j,xפDk��[0"O@��k��>�H��͐)�F�	�"O� H���KŠ2��e� �'��'��)�'aM�}�&�AB�U�䡃�v<��'�J��жLW�11dH��'���*��@�j5��Pj^�i��'m�u)$f�M���aq��Mo&]�	�'4����g�=_.��Ȁ =jB�y	�'�&QY�.9~���Z�F�n3	�'3p��#��,&�b��@�ǆ=�0}�	��� ڝ���ܫP��RV��t�Bț�"OR��7�͹G����LK�w&�}	"O�H��D�7XB��KI_66$k�"O���C�;I�����	�h0��$"O���`�2'r�"�nF97(bh�`"O��`Z�jk@)Aȇ�G"��z�"ON�Sk�%p(i���{\�I%"O�j4�&?C,eТ�-0�"O���5FJ��P�f '>��@�"On��E�D��B�E��)�"q��'���@ܬp2(��E0	f�)AP��<��n -AC��i���xU����؄ȓW�z��!(|=��Pn�(��*�r���b��%(,���	=]�E��v�6 ���>]lDXڰ�X-XTy�ȓA*�[sT�Fe��ZE�AI/<�ȓP��r�H�O������	t�d�ȓq=�}qn�(T�0��S
�N ��9=��J�Fڈ[ԍ���^�u��M��]�5�:>��T��;O-(���%;��s�
?&�'P=q�bd�ȓI�}���#���5 �"4�����rq]����y�h��bs`��ȓ��9r�&σ}��h��e�:8G��ȓ1|��w[���ڵ@��mG{B�'W?�;I
|��tB��F���b�:D�H��Z.�!�VBG*;�m�e�=D��b����HzF����y@@�l1D�p�1HYcl�A�d�*h���Ua�O����OB��*X� �BĻYw&����֚;�!�D�=:H��-���CcnK.�!��������^�g�ԁ`P.^�q��I�`�?E�DN&T��	9��D��� �'u�<���ο.dz��Έ:�)P,]v�<���H}â]:U��P>hEY�'�sy��I�\�<9 �G�n��l
��)Z��# 矨�'+�y?O��$�'nL�9��ǱWAR<i�"O�`���I>��t�  y X͂6"O�M���A�F�paIY�[��@�p�'��@�)�''[fi+t�?/k�$�SC�@e0�Y�',�1���D�
�x�U疶6`��
�'_q:a6jX�ԣ��.���
�̘'28���(^fC�3� �"&|���)O��1�O�@h��ޤE�j��&�=_<A��	D�d��&��^yh��'���FhH(Q��3D��Z'�J���\{ΐ?����B4D��sW�S	<��)j���+�ɩl3D��p�났?��)�#	�l@���G�,D��(��W���)�#��.��i�`g(D�`┬Βf@�t�� �9\����2D�����vVAƣHR`�5�BB2�%�S�'LV�5�sbF,x^�exs�N�x
�`��`�x�´�Јu�}`� ݥ[��$�	s�'Y?�1���	5'�3gÜ�L�8�G$D�t[����4
����"D��{A��mr�!�WN�3J3�Q�g"<O#<y��D�~|"҄:#��!R�C�<au�3=�ČY�C�2R��j�g�V��hO�8
Ѓ�\�*t��㰅%'����qm�b�E�0	��<+�d�; �����A�|�ړ$R�Q��e�ӏMp(M�ȓH�b�"wA�0�� �Eوr� ��U�F��t	C�(�[��< �uF��'>�Фe��R�����͓$!�=q�L2D�� >����G�$ReXa����:����O<��I��^���	�}���6��Z!�D�	M�.)p����Ƽ�����3Y!�Ċ?p�yI�	�+�&� n�!���Ib���4�X��{r��,�!�dW�"���1U�j�b�� H!��C�{1Hh2�\�6��K�*/4!��%Mrm��љ?9��0�.,!�ZhsP8���̝?ؘ�5�8@ !�D��kp`��r��[P�kC�-n!�DK�{T0�EE5C��Z���o!�ۜ'��ɚ'�.�0���O\!�D�o"�S�Ƀ*.{���.J�b�!�dž[=ލ�pMю\[�)#�m �&!�J$�T]�DҚOA�2�Jښtџ����C~�O��+�S�!�� ;�+�R����'/�tHÂ�w�P��U�?J$MP/O�O�����v��=i�ɜ&0l��@��!��#����f)�+j�A�Sf�r�!�$F�>���v���ayi#�T(�!��_P�-��=-V�Q����!���
N���٤iU�i��D��"�} !��=�(�Ҧ��	|@9xA��!�$&#A&!@�数qh�0 ���T�!�dH%+t��b5)T?RgR�A�I�!�d�ek��'�n-��R�g9O�!��%PY�)�R邳���'48!�D�����S'.�\�Τ��?2!��M}4��u@H��̛���!�$��r���)v�V0��t�!�Dۑ,���v�ԹJ���HX({!�d�q�x񳴧��<H
�j�׍6 !��p)QT䍬8;���g�PF!�U,ZG ]+���"L���1>G!�D�)_��[�%o

Tj4$�)!���&�h�%���EC�6w#!�dG�.j�Y(��Ԓ�������{B�G�/]���ê�=/X�J����J�!��)q\��`I Ha{��<\�!��W0
xP���T9P��5�ǃ;w!��_g��i��ڈ���Z'��6k\!�P�n��Ea�)�=
�	���Q!�䂙)��L��A.s�0�5�3UF!�Ȅ%��d���[�C�>J�F\�7!�$R�$�@���Lc�t�&��k�!��B
}�x$�&dZI��A�M)"�!�Ы?����J�G��H�b��D�!��M're꣥�N�hf
C�<�!�$A3=Zb��啍%�L�Q�'+}��)�'-`ӀA;K�$d�4�]���	�'��%��@�x�B�êYg!(�a	�'�r`a���i�X��*Ěr̚��'Zl����19�ЉQ$3s7b�R
�'��PYT�O�G�\;�O��;qެ(�'�����*X<�p)���9@H|��'����e�_$uY���O$I�n�����hO?�: h&&P�y�����[?~M:�Rk�<Ԇ^��<�c�`�#�	��
L�<iP�#dݚ�C��> �eaC�XJ�<�g�".����U��{�0����~�<��P�Q�`�LқFvD!2��|�<a���r8J�	*�"N��3��m�<	 Nd�`�Btf��,���{r�jx���'�d����Q�\����`�C��x9��� �Y�
-7Œ��"��TX�"O"�z�Ê�-��nR����"O����f��U)!n�̦�@"OB�� ��x�ę!�=�b"O��0�˄4��<���5R��<��"O��q�M23����/ؖ?�.�Ha"Oz�sɑ�k�f�'��g5��w"O<[ԓ:�l[���t��"O� ��KR%o)8�{��[kV\��"O�iqG���x֩)��[l9
E"O� �E��	H�u���V� C�Q"O6)����3�� ��dߕd�(t"O�P0�?N&@bd�����U"OdhA��%�r� V#�.���"O(�H��9=�N�����'Mr�8�"O��@#ǂ$�>=Q��i�"O%�c����ש�y �,�7"OR��&*`�,e��钺_�d�r"OlPS%�4l9b�腨�[y�<k6"O,ZG��(62��f�7ql��"O��i�+��͙r@��
r�D3t�'�!�� P�#ߌ�.�!P%���!�_�<�8��ŕ�r����S$!�W#`��Z�kJjA���Ƌ�/!!�*5F9��HU ~'b8y��/ !�PUl����+P��xB���\!��/aW�q ��C(#��-�!�$ŧgQ�dW%@Y���g�'y!�d�2H�D;��=x<!��e �`!�Z`����No΁�7��B�!�-KDB��B4e�lXJ��	�!�d*mH@��ƅ�"�xk�Iػ5!���n��]f���-`�J [�!�䑑-BP�A�-�D�Ca�ȓL!�d�5��Y�W�� :�j4c0ɘ�VU!��J6�8�Q0�YZV��GR� G!��*���ք�E��&��K3!��=�xq8����m�X��CőC-!��3J�6�5�.z�P522�Y�!����˵M��E�\X�F"ۖ9�!� �&L[�*��+���2���B�!�$Zn�� ���riZ]��˝��!�
_���X������!�!��ܳ(��ab)Z<W�58��Q)]�!����i�C��uX�e�<s!��[���3��׷ d�R�#łD!򤝛^UiL�&k�%�$"�#B!�DԆn�"��KV�:0˶e�0,�O6��Ӎb<pa��BtHe����8O|!�.]ep��^{�ݡ� �(I!��@t��� -�C����	�� >!�d	�E�.��Ađ gX}�D�9#!�@�e�����rZѻ1���r!�d�||d���%��`J82���q�!��aC��"qj��{?r�ʃha!��Ь]�r��X �Zt@ �rT!��T�B�V`p�N܄��x�P �"s!��a�IZf�ۿU�ѩ���2^n!�䎂f����\�0=�L��-�s�!�d�;ШT(Q�Z�̰
��p!�ă�9��ĺ�(ʅL���Kd*Ǭh#!�đ�J��|`'`�~���1��UB!��5HM�5�D��4\R��P*�!�D�2�|�1D�_-���Ӡ���!�� �q��G�$�^�⏛��FT�"O��tc��{���� ˹Ix���f"O>���Õ�0R�Y2�R7nB%q"O�X�a��� �V%~�1f"O����/a�0J�͓ x�xi�"O�Xd�߽o�V�y���ĈAxP"O�R�o^g��r��L�l��"O~�g��&B�u��ƒN� ,�E"O�x��j>A�6��d�?e�,ҡ"O������m�р���`=��"O�xE�N/��� �.Ӻ�[�"O�U�#��}?t���Ɍ;�P���"O|`aY9�����HS�,xe"O��8�!ڜXQ���\���jq"O^��Q?R��(qC�)@���"O�M�eMP�g���,�+�H��"O���� �z����R���b��("D"OH9���L-Lv�I+hS,r�r�"OJ�� -W0U� �'O[{��:�*O�<�AA������ڸI���(�' �4�1��.{
�AFe\+��Ց�'t�<B� �~:��f��%�}��'�b��'6��$as�� ���q�'��M ���_� <��@�TP���'�Ri2/��8V�*vLO]�.�c�'6���
�K�0�� iE����'m�aa!��?)n��m).�2Y	�'����J�d�LeZuǾry��'jB��!�a`d<�S���i���
�'G<UkA�'t9Q���e�pu��'LZ���o��^Xt��!�W�$��'9T�c�O�S8�;$"�z:Ĉ��'nyc�`(
�Bs�Yp���A�'�LdC�O>4�D|y��f����'ƕ���B�	����Dȉ�Y�x��'�-``�I�@���ÇU0O�����'�(���.[�Y�ŅFv@��	�'�@���E�o�b�p2�ܧ:�xQ	�'p�q��#Z�,��x%�7fv6��	�'�.����^�����@,��s	�'4��!��<:d�� l��1�e	�'=@�J��C&�D�a�I� C6ƍ"�'��!��'yĨ��nV�:�\X�
�'�&���g�*l�'�*+E��	�'|���?S�V5jb�˗"�Ri�	�'Y����t�q�*Xjl<�`KXN�<!�Kΰ9r��nN�dL�u�N�F�<1��5Z�L�)��0�VLs��NA�<�Å�$:�by�2��CB4]Pa�z�<!"�R���x���^$@Qx�t�<���79n��y�(��CY8}��JSq�<�FZK�<�s�JO(^���k��q�<�tI�?OHZ���h�V��l�<A%A�$�D��eb�6K	�Z2/P�<�B_4t����n�^�yrIr�<��ĩV:�0��E�h�j���j�<)�F�PJ����҈{�nL���f�<I�a^�[qh��S�s�M(TlWx�<�R��3��eX��/-&0H�lJ�<QS�2"����Ņ��h��"I�<a`��W�!��J۰b����E�{�<����n�D�2��0��l;d�z�<9�]�,2�hRg̨L���JG[�<�v!7
��#�J*&$բ��Pn�<� 4������(l��f旳0PN� "Ov���nRl
����_�R&���"O�;SC�B�]���� �LS�"OBH��j��^&0{��n�$1r"O*�㧯.Q�ɨ4�ŵ.Қ�81"O�Qs�$G�.�|�R$�%X����bǤ�E#ԓ|i�p��(g����E�Y�&����&4��l�ȓ\���,	-h0�P�ύ!B��ȓ<u�a����qT�1PqZх�2:�5��pl0�W���7�����y@��ᓅ�(8i�UZ��	� ��eJ�i��+�nG�Rv�^�g�Ňȓz�\hقCD�o��5�ـM,b|�ȓK�F�Ĉ�ۂw�ʿ�@�ȓo�ЙPOI&�����^9`���ȓC+4AE��Kw<eHݳ�>�ȓ%T
��*U�K�|��dQ6;�x�ȓ^����sBA5�~�k�ˊ�u{ԅȓ3M���1��RA6���$�#�Hh�ȓ.�>����e��9�(ʼ���g�,�T&S�숑"�1A�T���_�"L(�����-)lC^ڐ��ȓb�t�sI�5J�dՐ�.C]�ȓ|��q�g�fa7d�)��\��n�@�<��GC�0� �!I�e���(7F�S�<Yר�z�t�a�N<pbO�j�<����=$Զ�فI�;d`��Ac�<Q OШ.Ʈ\Ö�'���� �[�<�o�N����eW4XC�/�N�<�	��bt�� 7��>7tބs1�\I�<)��K�a���d�$�b4k `F�<�1J�B:��TK�A��T��	@�<�pOԄ��lz6�	`������|�<�.֜G��h�l^ ��xxv�y�<��nY�¶����Ϳl�N���i�r�<�@��A�`!��!�����\p�<)�B��CT|p�0	_�� q��m�<�����`�R�FD�M�0��_�<�@$ÁvXeu��r��Z��Z�<铨<Q��B�-ȃ �0��"a\^�<��$�=�p�ɐ̑�p삽�QS]�<�(	�?"Ġ��M� 2<��Da�\�<ɖ�ۥf; �#`D�n�^XQD�q�<`��7W^�()��T�l�
Y�1FAo�<)��BkV�9��M!BWq@%�^_�<!#�ξB�fh�gȋ�Ƃ��X�<9g���C�|1yA�L����S�<�	L�o����@)�[�����*�i�<aa�jd�l�Fngqn%c�Xa�<�c��7�H]�!'�*lL�H�.�U�<a�@��{%ب�w�(�8�3�F�<�b �Y��t��@(wJ�p)2�M�<��FYC
��ا^�0���b�<�!ND2B��պ�aW
-����Ɨu�<�Bg��!��z&,��x��l�<a��Ӛx^� ���tj�XfbJ�<���9M�-(��܁tΘ�@�I\@�<��	�=W����WF�DT4��Fz�<�f�qX��P iL
9�4�l�u�<�R<+��r��f��t��aIj�<�c
�
}�5d.ڏm�f"!hI��<��g+��+g�Pu��0��مȓ^�P5��0m:R� �)@0SI2q��S�? �љ��2]h����n��˳"O`<���S�X<���"��!ct"O��p��!��q��C�-�"O"8�dk |o`˂L�&Bġ"Od]1��ZbH��*��tn����"O(l�W��L���P)\xP��w"OP�j%,�N�0��'2jy��"O&���Lp��q���4���"O��`�f�$�j��ƍ�,��)3�"OdQa���)�T W��0�.]��"O��Ȅh�5q��=ׁG:B�0\{�"O��Qt� ":&�u!G�4�N�"Ob�hEz2|��Ƣ�F��i�U"O6ᒂ$_�	��p�g���/����"O ��G�w+4�9!k�8B�X��"O<���W�H9H$�%�[s�3�"O�ha��A�1(�QR(��4��"OH!Q� �	Up��gF�<%V�UCt"Of�뢈�2��y%	wF���"O�`͒*H�I�W��6?|t�#"O�@xs��h�BP� ����"O�ahi���M�6�i�2��a"O��ؖ��m��#�c���s$"O�L:ؘ9N���#��|�1#��!D���p	�v��A�C�#��]��',D�ru*x� �L30Z�mz �)D�H;�D��1��HڦL�~���	�()D�L#���8r7�Is ���%�(D���v��20�a��#�hr�)�5�#D�Ԉ��J>\�JtB��et65k��#D�px�DA1jC������1Fb���"D�D��a!�ى�hP�R����$D�$�G��s�d|�@<#OH0��� D�$������V��֡��z�,���?D��7iP�g���I���"t1D����d��W���Q���Zԉ:��"D�,�`͛�&u��Ibc��!��`�v&?D��@#���*G�-c5�.Q�`��j)D�t�a�m	:yXw��[�� �F�&D���� �x4,03��P�QUڹ�&�7D�t���<.�\�uH��:R�<I��"D��1(D�{�x"���)u�T09�d%D��`d��cN,%A * +ьd�1�$D��Z�j��Y$0MH��	DFx�%�"D��j��p9��ZGDωkIb@Q�?D������Pn�](:(Y0�!D�К��"�Tٳ�jɫ:��Q��>D�@!�)>����F�7��<D���uCZ?~+z�k���Q���i�e5D��Ԅ���t{ �'Mw�U� (4D�ܱ�[�_��Q�#��R����E0�C�ɞ;و�2�F���fȒfs�B�	)��}y!@RQ����э�=N�C䉚V��|a%H��p���CdN�3�OP���B�U��Y!�g�UG\�0�FS)�!��2?	j����WNn��T�HNQ!�$�F,pö��8oJ�`���C3!�Q�S�*�Z��Jm�Ux�P�~�' T}��	%�^IA�Z5P@���
��z����v�dX��4r$@a�@��b�A��1D��{�`à�4��pA�#���k,}�U�<�O�"<A�l�/ �e9�ܮ"Fn�yB�V�<�6'͡ts����!�.C����5%j�<��f�B�V��H�Y��2�$�O�'-Bi�V�π 2�� ��@�"X�I;d}ڣ"O��R.�_�Dk��å	v$�ē>�'{�O�|P���K� }���C��V�"w"O.�Ht�R�G�vi��Q>!v�*��d���0=�a�T-s�:��Q��6"6+A�y/B O�1��)�.%:�������~2�)�'S��!t
�jŰ�8r��<b��?QM<�Ba?��4^��*� ��;��[bD͔p*�C��&4�z�8����Ʃ˜.��=�Óx4�y�5`ŔZp�9k撼na�����D���`_��T�M�8�B �>�#�!<OTH��M�7
L[t�՛o�n�kF�'ў��$_�%�H9z�-O�">p{�f/D���	�2	#����Δi%XaC )?������'�i%-� ��)����*@((�'r6 ���0w��яX,Ib
�'�,���(��kI�4Fj.A�'i
�4�ܮ/"f���e��>-4Ũ�B�)�t ˀ=�,��ud�Vⲽ���)�y�'��R{Ĝ*�*H�K�4%���hO���dK��xɖ�մX~`�A`�F6DP�W��(��Y9�'����19�EZ�bF�L��']!�DV!�(�h���%kHؽ� MV�d��'1����=��ڍWSLXS'@;W�D)��^o؞�=q�LJUÔ0ٰ�߄[D��H���g�<9d"R5y�4Pe�G$�X��Ha쓜hO�O ����F=I-2Л��O� Ȅ�;�'0h��O({BM耥ԎpL�u��dCV�4��ʲAI`c��ԯb՘!�c�$D��і��*Wf8B����`�أ�x����$�͟T����$�� ���BE�#E�7lO��y���=y&i�.�TIēr�'�m<h�}B�d��dղAڶ��5���%�NN��>�S��oQ���F�dl��#
%�)Fxr�)*�틋K	P�3��d.����Y[ܓ��'EQ���-]�xeb��^�U������n������[n�4Ц���]�xd�����c�e��I_}2���Je�W��Yq��� �7�yB��X�=�NF�`�Qp�L^�y��IP��g�8Y��r4�ȊE�����)CC��^��\����5"�����A��ʓR�IY���I��
ﾁ@G."}��EJ����#K�}b&�|}��Q-&���x�d+@q�N��y㈎Fj�a���V�0H{�f��?I�'�����W�w�r��2�|��	������+Ч�'�*=��<a��-:v�:D�|�7��$*����ް#MxlL+�	��$Er�O"���-���2�$��_��J�yb�)�S��)b����K�D��$OT	 �n��hO>�Bߦ\#�=�4*Ek}dE1#��<A���I�h9��W�`��YjdK�<�(O8���Vc��RK=[!&�+t�P�=�a|��|�k�:L��aH���5�@�q�^�O\�=�OPF��%.��(��#6����(d�'���#n�^H����ˊA쉡�'*���
�6$)P�ХP�)�{b����O6�t�R����2A�p	�`8O����v��o��b☙j��ǍGL$�l@�<b��E{��t&^���
�����0&υ�yrV�J3<��"��жt8� ����(�O�9�� L�`�"2���s�^EC"O�|2ƄsIU�EZ=��5��I��y���OT���`���fN�%����"O��xAO-[�y[�O�,X�Ľ��"O� @��aNդK�^�B9[}���c"O������ �\JC��_hR��#"O&���.�05�h������ک�Q"Oj)�7J�+k�� 8��L��6
��a�O%j�8�	W�#g��pi �(쳎yRK[���O��|����44��p��O�̵r	�'x��JB�H6�]����5>����w�)��<��J\I�H�e�P4���	%(�b��}؞,�0�^	4��вe�,wJ����F_�.-���	M?�PM^US2��R˺@1�8#�����hO1�:�O`��`��P����ϘYłL+4�	��]mZ}������[� ���o�iz���H�:�y&+��8�� ]�4�Ќݫ�����d�\"~����"%��2F�Zx����JG{�'�ay2��6�bEַ��Bb ���xB�U�PVa� q���q�H�{^���'x ���Q�&�hGɼ/�1jד5)tc�rUGԚ&�:�����zp�鈕�/D�,�G�lnX��R&�^کx�,�	Φ%Ex�x#6>�z��i|D{�c��'^#=%?�{��e��\�@���rX���n'D�� 0�G����#b��qo";wF"����'I�<�1D1|@�DpPb�P.�F'
w�<�W�#�D�� ��AR�£%�q�<��lϋUu��8�L	G(Ų��k�<�%��bER��ł?`�c��l�<1��8�vl��R;�;��Zh�<c-�yc�!p�È�I]`=���|�<I���$����7B�M��%{$z�	g���O�2$Ԏ��ېt��H�[9U��'"�ce��l0[��C�W�t��}�'�LR��@�ir�P�����J�ڵ��'{N)2�n�F������ʾQ�|�
�'7�	:��o���T��;r��J
Ó�hOfhXD�ˊ&���A@��Bx@�3"O,���϶b�1󕩉�*� j"O�{	��[����åSCk`�3�"O�[��k�Th��+y��%;`"O2,�tI j�j�թL1c}I�"O`(�D����t���Ά*Lr(0�"O�	��Ђeb�H�f�Z�\��"OR q#"�����G�I��h��"O��	�j�"|�J}���d��lA�"O�i�(M�>-1�J_�+Ԧ��"O����C]�3���*M	��PS#"O�]��-R�gЀJ%[N%��"O�<�"��Sٴ%{Vb�1.p�@"O�H�1b��D��q���J:ThH�U"O8̐�D�'E�\�����~���;�"O�"�5��̳g&�(��)R"O�3t�_�������G:�j�E"O���a�ӹo�1Ö�pĘ��"O�Ī�U�6\!�T!W?��Pr"O�A�SkZ���S���;���y��{P�DA.� �p�%)dy�ȓm9�=���KFJ<ٶ�Ay���ȓ��d��Z�v)揓<5Cm�����B��!}NT�7�<0C<�ȓ!�mPV[HTX��O m�v���Ir��E����u�F�@,�ȓ_�NmKdmK�0^��J���UwQ��Q ��RF��\d�f�γJVڬ�ȓ:^2	e��u�D���3��(�ȓ}6��DS1A)Ĥ��!��̇�S�? H�z4`��lR�pA�T8Y���A�"O:Y�	_/#�ʕ���+{Kp"O����>L~���<G(�@"Oq���:�����%Ψ�Z�q"O��	0@�"<�4t�c#�Z���k"O��c��3��h²H�6����`"O�-0� .����&]�>�D0��"O��I#�2�uph�
5I�g"O��a���MX�Ų��M
8����"O*�$��V����h��)�u��"OH�#�8���B�FE���0�"O��#�	�a
�D�Lt���"O���5%��V��}0�S-�E �"Oε{p�< ����	ӸN�~pQ"O��i���22���WiZ�%�y��"O� 7^�L�<���	�&$��"Ovِ��F�D1�d插F�>%
f"O��Mȸw J ��e�7u����'�N�9�/�,o��� ���N���re�+����'/Tt��D�s���`�'XԠ �'��d� E�F�Mb�'��!��'$2\;��
?y6B��"]ےa��'�~Eh����<��A8B�p�'���&��k��,�����ݮ���'�����ґK�&�����"��Y�'���Z�lZ�r|+�&�j�����'XT��F�ի ���Z�Z��'K4Y��<j���7쟉[��=��'�"DP�g���*��R�Hh��y�'�ҸSf��8֌p�Q7Q���	�'�\9������lx���S�\�@��'���{d��pr����`�=O�l�P�'^ ��Ö"a���'�*EMB���'>D@��K�7� �x��P�3�u �'D`���,��,i���S�*QA��'+T�jR�4"$P�%8 �����'ߘ�E���Y��u��?�P!��'U�T�0�[�0�I%Ɍ"A=10�'���J�^�l}
j�i�|�	�'&ZX�l�)��HHwaB�W ���'�؀ǄO��t�!4���'`���uA�,I~�`k�I�.�y�'���h��ϱ��!�tc���� 
�'�Lm�g)ڰ����T/̕i���(
�'���as���_N�Iy4��1)�n�h	�'�(ě���8s���V�@
#��Q*�'(0�R�)�z�2�i�����'�u���ox�T����as�'��ᣃ�n�L���N�:cV�d8�'<����eS=hr�b�!H�d&TQ�'��3��
�+�\Z�������
�'���5h�yB2�I��\�	Fm!
�'���!��/��" �?~?��'��)Qć]�t�8#�m*���'�4�CR X�R�y�m
�c�"���'����I��P�Bw��A8�:�'Y�J
�s�j��f@H�8a����'��L0�\��&�ތ*��a"�'3���=I�HA�����&?>;	��a%b�12%^O�:�q�HCg��� �� 
O@���2Ct-��m!�a�LQ�D�D]0Gp)�~�5(��{�,	�1Δ*`�Pe�AL�<��h+�ەe�$8�D������<���I1^^Q�#j$}��)�	�|�� hG�E����E�/(!�� �Lb�@�5?n�xeɕ�T������"��)9�"%�'_6-�p��q>a
Ԫ��왲	��B�r�J\�u;Bo,/������=1Enm��?�PYB�/w�XA3Ca����?�+N����b��(mb�>ыa��$t�+���1}d�]�@�9D���<�V���Q�*@�!0r�v���S/����"�>E�$ofg&ت�I��3��p�'�_��y"�B�R��]YV��-�lCwH����P�P8��&Z��p<yL�$ᓧ��}�Xa�c���t��8f�����PѴd��	���=;4�?)���&�*���A	xD3r�T� o��c�D��,��	(v)�nPeX��ϵDY!��Y�9�)ۅ��{iHt�$�1o6��2_�d$��&d1�O�zkL�Oju�q� �OcNջ� X�4�|�*E"OT�Su�̣{c8#1�M%3����>	f�\Jf����#���Hc��1��"��Pi��	��i`#�7YΔU[�'�$L�C��`�ڀ�ԏ�,F�@|J%&�%�-(ބ�O�lS�����ē��Z�gE���@����<��-�ēy�4�YuH�#��3'��F�L�Ӵ�S�P��\ �n9�O���h�+*��t 4E�Hj4`��'Vʹ���*�ܔ'D:� A=i�4��ď�+Iإ 	�'Ȧk��7#��ź��=)�h�CL<�%��9|]0���H9��^�)a��J,HT0�Eeǉr<� ��FL8a
�ݟ_������`5�qddS���	1�~؃��L<���9���Y�	��vQ =��ZH<]�J��S0���aK�GЈ�d٭B�$-{@�<�O��X��X�H3�,[ďI�_���'�l(	v�8��9j�i<�᥊X� �f�r�� :��sr D��DPҽpQ��P$~��' ��M�\��e�N@֔�Ё�:��O�bT��Ą8a�H1B��R"%������i�f\�p�J�e�L���`φ_J��Aa�g���I�l�k	�t�х��J�AV�*�3�ĉ�K�n�b��=<\�D�#� T)��X�6kȕy����|���%L�t�b��!�J͂5���K�E�d�7/�<����.[����| �Q���ӳm̘�q3`$t��R%��q[����>5���ٙ7�]ay���r�K56t\�2���+�H���BhH<1үٚ�$pi�g
�"�h�pD��sMz��a�
#C�;���-H��'��X7\�zt�̹+&.J�(P�;�~�B�Nx����*&D
��Ԁ>/���m'ٶ���"C�v�X�Ӓ>���I�M���
�L�=T	�ið'K�>�>������<�{��>�Ӡ
�<]#�J.��s��s� ˓6.&�pv��4_R���䗨^4�3�a��e�N� ���]�$�!L��G���)��K�J1��*�+�(i(���!A	�� @�	:.&���'��i����	W*$@k���" �U�J�@���\QOP̋$�3O[�m�j%�4���(4�+tu@�c+<���J�'�V��#C	! @��`�窩p�*Ҿ{CʴB@BB�RP�P��J�S�O,Bha�I֟G�&��С�!�x쩌�d��N��(�!%�S?-cX 86�ޞ`T�=y��=A�C�I�N����7B��i�@��3�˱Y��ʓ	����.�)ʧ?��N��8�)Fj\9f��i��?� YQbM�h���)�^6l�Q��<'zzӇ	n�h�0-ѫW�8���C�R"���dmP�1C>"֑!$j� #X|�Q�V��Hg�O����3N�2-��j��ѡ2$�-;��.lO�0&ļgP�I�7#�)s�́V>�@��f�"? hs�O0S���I,bݘ�+u鐋mnҐZ�$�X �*��ɼS���%��Rp�V�oM�d��74nF1q�L�?���d���<R�J� �f
!�$K�{�"��kW&"Ԍ9�G_�|��=�|qBm�{�1p��ź�`���X;�OdͻW�Lx��4r�(Q�	74�ل�I�/�m{sЌV��KM3�Z݁ !�2$W�4��A@����i�,<S��o
<Q���B#=9ǁܙ$�����b�D� �@��ah�Q���0M�����Ƶj��*�N4\�Q ��3kX6uzրR�-�(!3�������@	,���C�<-����*�DL��XT@;/9���ɱ|��ր�*3-��{��`#�̞*.]9������D�̞b��a���U�cVB��7� ��Fpƶ��D�!�= �
8n�	i�̛��TLY��� 6�$����Ywμ��� ��N2� d93����y�5�歐�T,��Z��'� BX�p�n1o�M5^���"����2�@�(k\d��պz+.�)Y)����&��M7T���4A41#s%Ё]T��I�BW�d*�jĎ%0n�
p�\�>],�	��B�H3O���S�ÆG_�t:�O1j�" 	\�<Y$T0D�?�ժBmɻ*[t9!	�3fpM��,(В�o�.f&(�HV#̯*%v�G|b�^Ѽ���ϐ�F�(�Ԏ�Iĺ��e-�K�]B䎀�L�>\�4�ˏ\Զ���P%E��S$a^d��w�F�K|�@BD��g��qj�O�x=z���'H@X��_��v��� a��80��G�%��|S4��:S{� OB�|pi���7E�����4U��C��<6��V�ʡ�EM5�d�x7��+�HOZy���ũ\�����'3T��S���?�2�옫rL���c��;y"��DM?˂����>��#�*~D���'��x0d���A�?O�0ق�� 1V����C1�,xYR�iYz�@�F�>^|Jy��.O`�I�E˺�"�U�QP�J�_h�p�5�U�W� ��Qb�W � �N�9YLXM�'� ���u������	v`d�	��P'a���RK�;=�$�Ig��SN
aJ�K�<,�v��#K��skr�A��f����"�����G\���S!v�L�#n9W��HU�92� 
�s�&	kP*��%v�5˰B�cu�9q ��>�N��o^�	#:�6���l�q�3o��$���

��A7$�ئ��'R��0��v���HH�4mk�-p�'���OD
=N�nڔJ� ]Smޱ�੠6���N)B��".�>~|z���,hD|؋Tb�*�F}	�$f
6Ċ.O��;��D���!��'ծ|둪�3M�<%���>W͚�h�4o?X�C��&&3\7�2% Bi�RM�w�0��dG)#�JRbT6.�j����	h\Ez!��v:y�e/�o�ޝ�'�(|�P�� yޑ� �rK�Z z	�c/3|<�,G]�/�\���bW9�-ˇ�#Uz�1���Ś_*h�s�2~>��	}�}�FÌ�{u�)�\���[��&�O�%�P��f��9@Ў'mN 
WHT=b_Ass'�,�X�� p�@�ƅ�45r�d�P�#gZ(J7����+,O�,�VE��}�+��GL�mXqDG7��=q�d^@zl��Gi�V�k�Ր"�*1��G.@~"Rh�>G�Vib��!htP�BD!Ǡ#�T�?���K�vN���$
h(} ��W`�'p�"�MÖ7�%�L�� ��E�.`Y�L��Ip �q�	�n��Je��S�쥋�'`���V�NUO�m�+ʾD�����H9ow��X�'P�)�%D'4M�Q�3gǫ%�2馟'��3J�n�cc�G����6Ұ�y��śjl�X��M�7�`�2�,� N	T����I���XSm�����Y��x��'w�����Ξ_,�-�E+D���Ԍ�e�h�̯$U���fӘ�X�Q?Pj�ѥB$���d��	�&��r-Z�on.�)≞,9�{�Ƃ#������M�ȭ�2煅13vA7��Q�985��JH<�V-�^��9�ɚ��*�eU]�'XR��fMw!才Q�Oa~�I�b�y�T5�u���S���;�'t��BC��)¶yP�jE�T��1s��4u��2L;�)�'4D��a������Y�EP O��1
�'�N8����=������r�n�{	�'4(�؄�є��\ՁZ�fPh���',KňWL�t�Z�nאhPT ��'hH8�tB޹!dy��VS�:���'�P�W�ݚ��y��a�$���X�'����6!u4Ekg�����(:�'\P`Y��&AL:@��(ӏh�
�'뎉 �R���zt�ڥF.�8�'����兤J��Hc";d0�3�'�n��OM�E�l3B��=yY�'*������e�	t\�����y��5=vh������(��ቌ�y�Ɗ�}I��� a8�� H)�y�ϏV.��e`@	{���X�͝��y��S� E2OƁpp��EC��yR.[:�,d#�M��r��})�]%�y"�>w0ܢ��B�v��[
��y�m�6d��I򱡅)�a�K��yI�<������)�����`�y�G*~,A3jל/j����3�y�I��%�i�A�RcZ��dԕ�y����޵��/_�H#��zT��y�H�
=���Ca)�
@�+�y�2n�^���l��8�qQ�@�y� V-`��-�#�[7('HH��"E�yR�M�V�h��4L�)}��3�ϋ$�y�%�:_4@e�`�-~Bqpt�
�y�� �V�CCU����t��y
� }�ň��rE��G�)��Q"O A`���X�!`�@�T��T"OR0�A�ܶ �zD� �>)��(��"O��c������ToČ``m��"O��������)b�Β?��eKG"O������$���Ć�� q6"O�9	Ԥ�6�^ ���P�i��R�"O~�x��е	�fP��ՐUG"�"OL��2'Q�b�n���k pԳ�"O��jRo�rXF��EE�\ ����"O���4���zd�3	��LN� k�"O:ɷ���u����&���"O�����U:?S�Pt�[����:�"OXDbe+@�$lh�׬^)TXN���"O�$��-��p �"�U�Y3``�"O���^�;<d�aM�I�+e"O�MZ���c��$B`틐8�X[�"O\�{v,[�*�b�&J,8�&�0B"O�-�����~O�����B���"O�i�E�,�4DX�ē�b���C"O�� �+��`��b�B�*:5ra"O�=+��F�.L�k�e��"O6yע��Lejq�U� ����"Ot�
Vb�$8v���	�r�8W"OĠ�0�O�Yf�X�A���Q"Od����Ar�сU�P�S�M��"O�ɴ$O 6y�ё ���.�  �"O�)G:bg�A&�6lrdXq"O$��N��sI�MY��X�{X9��"O��Z�"����Ce�4W1��r"ONóbʟqG�y��~�<���"O*�92��:n�!c��X�&�Jv"O�̙�%�J�ԙԇF�@8�%�f"O;R�N�(�b���MP�A�-�1"O�ܘv+��r��) �!E�A�*ձQ"OD`#����L�1� e�����"O(̸4�W�f��S�A!{��<�`"O�HB�}B0���3z��0r�"O���ܛr�r�'���,�( �"O�X).�4B����)	���q"O��� )Q�'�J�TA�8X��"O�\Hq�p�`�����C)z|rf"O:Q�p�2
���4��K=\`[�"Om��h�1H��T��9^+$ K�"O���w)_&	�  �,K�a��"O��Z�*h�!Pm��{)���"OnT)�mQ7TJ�=��S�4:|�"Ot���(Y�N�����eZ�R��(�"Op��"�S�_�l����!�Nd�E"O���儂���q@〱}��dZ�"O��r-IK@�o]�	�C��y�E���@� ��]daCL_1�y�GۏN:v$c��F:����N��y�@S{��rщ�sJ�)s�)���y/mi�}���P?h6��ED0�ybɑ�w���HC��#k ��`J���yr�� 1[�h�s��)�N��U/B;�y�I��wS�qR�W�?�p�$��y�f��dln���$�?{u
����[��yR�=3��hP��5w)p�� N��yR��'	��(�cM�y��˩o���"�N�3B���yI=�V�j�E�,)�d�I߯ݰ?�K(#x�!�@E�%rWP��x:��y��:4�� `"�Ė 6y��Y!?�飃�I&Mf�q!�w�'}��0;�
Ҙa��xa�o��xn���=z�H�7�B��Ȱ�L=��zA$l@�n�I��ҧ��d�adaոKn-����`n�t�S"O��2�&H�X<�x�P;AE2�3��p�����s��|�G�' ^$Bv�ڢ[��dB6����T��hb$Uc1��0n�[u$ 4%�N0[�a��#��Y�	0�42҅�$>�p}YG�
Qg�l�b	.�GC�x�4��,,���>	�7FV��f� �n)�2�K &B��!S�H��C߶$70����<���	�(=�]+�Cұ�S�Oפ�(�G�	|1�,S�F�����':���J;%�ʗ�?]:���O�-4�޽t�`��Wd^uի�;Vʘ-���
ن�I�r�x�B3ꚃjh��0q�Ю9@q���ٷ0�4$��
On,�E$7 �@*ίx�D���I�'T���D���"q��9�� w`�p�4�ʨ�����"O��%��1GV*q�QA̚z�r�'0O�[E�Τ�O��%/9.�%� ��)�)Y��@�6q�SJ-D�l�V�4*l��)Cb:Pܹ(}BƄ�w)&��#G^P�ɉv-,��cW?Y�g+�T���'�%>�8��i&�O4Š��ּ15���G�@|�4�	�#�Kl��(3<��	���`�!��x�K�	12���҃*)�	Cvn���x��f�D��fæF�LIHP� �X�:0!6Uni>d��I�V`R$qD�z�<�7� c�\���Ш���L?��D0I%�l2�[�`�\�&�
-j!��Յr��ܲ�KE�8��y�h,`�'s�)�3��;]ʴF�T!MX� `i$�����Β�y�I�,��5k��Kw:"���b�,
L�(࢞>1�IE_���'-BWc�x�	��(��7ܨi��'ȡ�"�B�Ĺ���3~\�RF�;e'��y�Kx�`�DA\(]8������K�AT��ay�cJ:4�(2'i�da\j�~�ؕ����lB�A��4(�B�I��b�{���/c�Ȁ)�n�F2hO
�1�`\(S�h�x�a�u
0����aθ0�j@����6ne�5����?i�!N�1;6���`R�;g��A�@�bټ�����i,=���9V@9�۟	94b>O�ع0� r_t	p���
�f1�a���x�����c�'y�B�@��ڼ �����cG�\����4�ԋV��0���[4b���>,O�A���R�l���f�A�XG��	��O@m�%`ĶP
0�2J����	o�|�U�ɜ%��qвl_{��|�1C[�A�r&#���}�ē%�s@m�tw��2Ŧ"ր��O�l����'A���  t����.}"7��!
u�[���c��+ ��er��'����F��.{����䇾Q���)�B4[W�!�7)N�_Gj�{�LOP*��h�~�(�Y�yR�))�%���A���3�s��M��E!_�b>���-��d�#� )��T��o�<�ӭԌa��p	*,O������~M���pD����O��T��s��3J���TDkݐ����� ?-�p� ҆[��Ri�N>��x�CT>z�b�ᬊ��,�z����w-dq�U.�d~���l��|�O^LQk d��|��\0#�&r��

��j��`	5MA�#4��(�pz�p�D�n�dL�b�1�����,�)ڧDv���&G9~�q2��0#�F~���7<���S���%����@�+iBH��&��!��g�6��ЎޟpF�U{�ā8`�	;{}��G�哒x�����:.����(T(�B�I$	Bp���z�hL�Ɗ��вB�I��=�`�ƫq�f�hGg
>l�vC�87�<�+""�%|�S�J @w:�c��û# �P*O������O2 (�!
!�T@��E\KB�'	�j�肃jH��݊{�@�$'g�ez�Ӑ;�ޥ���1yb��A��Ν��x��E^����jW#;Q��-�~bF�n�ԉs�Ȏ�?Uӳ���z&nDʶ�Ͽ��Y�-�h=�N�?dNd���)v�<��Hىc�V]��HD?��eiE .>���pj$z�L�K�ݔSJ��z%�'�擁V���4��x�D*c6¥b�e�z��{rc+u\���Ǭ�ަ9��jJ1�����ɑ6�|�P7&��.��(�p�
����W�vi*8�Ҋ�3�HO&M(���!Wc��P��4i&��՜%��e���ϊ�?!��S>�F�Q����� 8 *3c�1#�l����q�$ã7?�,c�kAFX����@,W���r�J��*�$	=|��I��?���P�E���G������K��:�di�A��ó+LHqv)"��Ak&D�@�Y7�L��b�YQ�r���2�Ak�E�/���ԫ���aL �g��C1���dB�iھ��{v@�x�t8K�ҔT��P@������=YUn��Б!  z�N��"g�)t�<�m�æq�Ɨ� Nx�s	ԻP�й����M�2�w�;�B7�8���)܆�~��˰�x%��
�$��Wlɮ�y�����T�~���J7�ʲ�|�S� ��,�n���T�:]�����ņ *�D�q'Ƶ;B%���
�M�0��k?�؀V��(�O(H��ϼp�n=�@Дl�ܥ����5[���;�ꖢhYɶ�ݚ�,L�'U�M;P��?��@�0v��Q����=�P���AW��@2g͟��2Շ�I�9�<M��>.��<!pFPG�6��e�	:��X�o�g Y�̓>Y�©�������CO�d�W�%q��l���J; wr���'4�������5G\Y�N��yrȓid�d�S�Ӕ �q��
����q�( |�{`��3���p��[±�r`�}y��l�I���R�Nn��%vk�dm��^���I���.M.�\1ѵ��`���-��K��5����vu���W`L%!	h�c��'S��y/O�0�K�n���qO씢g�U�~����_9N�ђ1�(yqR��'m��oL졛p�.5�Χ����d޻K��9��񉱎�O�n��@�* �#���ܙ��j�^X�"DeG5G7֥/��Œ���I0RR� ѐ�_1A�:QA�Y�J�$e���=s$��HS6�G� �JA�#$�<)M>}ܔ��}%fx
��%C�LXFzBB�	0��Y�oZ��q"�&E�XD*�&�z�4���aع)�~�����Sj򐁧B*,����n�OZ ��/}be=�S9R�ޕX��F=}��D����P8�6�];�ĐǏ�M�R���1�P�C"��E����-F�s��*vk�Ent�l�n��dk'@
/��n��l{ *�3�$Ҵ3�,��"�ߡF���$C(Qk�MÛ*���!L.rX��qBd�t�o�!bx�����y�)�b�P�Cc�D���f̖��0?9F]Lk+㏍;���j�K�J�$�� �5�ؐ#��C���T�i���'sў�:3��Zr qpҤ�t�"M�'|O��iG��Fr�2۴KB}B�-Ԇn�$���GM"T�dT'U�Fi��	�M� x;�� -�(z&�:�l"<I��ڌ�BI���)Q؜��	Z=Cl�}�4r�-��O�*��w�/��䈓�݂<��	�풊z�4��=E��d�P�0 ����eF)D�A#(D�ȥ�PL�d��CGÚad��Y'%3D��2��@�΄�vO�X��qe=D� 9c��T8왅$n�=5A$D���a�
0*���@��)�e�6�$D�`��˨z�xP���-�����y�(E�i|�yp��r�~��
͔�y��%>H�"U�Äj� `bsL�-�yB��Kp�@ƃX�X��͒�y��F�Bd��Iᣄ�'��J��y�d&~���E��n������ybϕ�ZD�v�ޒ	RT5r�@@�y�+�Q��T��_3q���Y�O��y�0k�ԙr�L�e���0��N��yA��x�N��F� QNz��M��y�g�"T���@Y��];f�ȇ� D�tO�9ؐ$r�\��j�X�2D��[��H�l�i3`��V�X�d�.D���'�jj�
�2g����0D�����&"��Y�'g^�D�Ųa`/D�0�4K�	�� �`K��C޲���K>D�$K��B�1ʹsT���h�8t:D����N�J#ƭ�-9Ulu�a6D��k��[�Gc���#X+~����u�6D�<Q��"��!f	HM��;d@2D�D�U��H� �#/�Iq���`2D�\���'-l�Z� 
�"6,��Ӎ/D��3��_;vQ��RW\0
���-D�K2�c�b��	ѾLZA���)D�$Sч����9{�OZ�T9bv�9D��C`��s�HL��� o����#D�P��A�~%t(�׍(��8��� D��Xe&\0hB��P?��l3q ?D���vO�6�f�n��y0�TS�=D�� �+����`��u���U�"OR�!�m�(-� �!�5>�<t)�"O�xHw�]�%�}�c��aK�!�a"Oʹ[�	��0�Ɍ9ԩ�D"O^�B�M/Op>��'�>p<��`�"O�]P�-�h�@�"�hJ�C:��u"O1�G#�0Z]2a�
\80T`�"O�Q��e����5��D~yh0"ObRpGבP� p�. 5,����"O��b���'])6�c���S1hЁ"O�]x�9M��t��Mů)W���"O��14��$V5��A�]�@��!"OD�XHJ4j!h� ��	|�h��"O^�{"k��c2n��K\�'X��"O Y	1J�_n�dj�*ӂ �b"O��S�Dhi�� z$�	�"Oؘ���J-/G��4��4cVER"O����"ܚa8p��'@ԥ4CXE�1"O��ɗ��Pr��2� 5��#1"O<ك���A9rY8�N�a��!�"OJUq��K���1Z��]�w"OhH�gk�8ZK��y�cU��D���"O�蘁ˁ�HH6��:�=@�"O��إn		g��9�K�J.�E��"O��R"��GC� Ò`Y�K���X�"O��	w��Z	Z���%
���U�'�����;tv`P�nD�WfZDœ�L��|��'m��%	X>yɄ��0D��'.�� VgC�8}+���"����'�VH��B�_��	�Z��'{ ��&�ĞAWty�U�F�(ި���'��Mr�!�<!�~�kei��$�,�Z�'~��!%� ,z�S�O���
�'�d*���,("t8e썉#��	;�'�<}� #�(4~8k�bΈ��$x�'�ݒ����6<n����o���'�eK`�Ő{�@a�En�=.���'"N�����;p�x��-�6�2���'X:U��D� �rD5�+��D��'�x�C���=F���$�,�(\J�'������$J�s��ܓ�8��'3��Y���Z���{EI��
=�	�'ovq"Ѓ�
@:�� J��/� P�yb�5�ŞK�� �)�#C�`�d�Ǐ'Ap��'��A��ԟ&I�I�PB�JWm��!�p̚�%-6���p�T���MS1���h���ݘ2 A����	
BDP�F�#2p�i`�e�0t�S}�O6�u;F��W�T��+[�&�b�q#�$S�`���~���y"g�f>}�T��:7�����Z�y�A3~2	S���*��,"1J�'�y�Lϖj_���&��\�`�ݎ�y���:$��Ή��у �2�y�T<P p  ��   �  S  �  i  h)  x4  f?  �J  %V  �a  �k  &t  {  I�  G�  ��  �  8�  z�  ��  ��  Z�  ��  �  k�  ��  9�  ��  �  Y�  ��  c�    a � � � ' �/ �5  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z�����W��K�L12$���SO�\1Yd�	�O�!�WR�H�Ī�.b�&hb1[��Q�|���T>�%		i�JI����z�`��6#1D��Sea�d]`b%�\th35D������?!�-Q�ė
?<��F.D�@3A�	5�Fy�B@WD&�H�!D�,s���CB>�rR�>dwA�*D�$0R�Ō*���B��30�)�-&D� c3�jFM �jp����('�ب�^��*�\�Xi��tU<Z "OlA�g`�$`&�@��I�kHH\C#�'ў�
Q�� P���]>�h���$D�\��.�h���p h�X�\�L-D������~`&A��K 1.V���5D�x�`ך_s��:��Yd8�4?ю��S7\�^5 A�ݯ�R=8�'��B�IP�&D���� �DU� �#$��B�I*1	@��G���J$E��LOO�JC�ɨp�\Dhfe�?`��鱺@�e��=O��i��b�x�Y�)[�ks$�ȓk��b#͔)rNQ��K�j>-����@�w�B�[*�� G<@�-�����DNA�R}�U�$���g\�܇��i��T}���.Ƞ��ĩ�C�(��C�	\?ы��?vԠ�F��K�#=���T?t���N�\Ry��:D��ۢ�b0t1��,�'b�tg8D����d�M{��CK,h�����5D�g�7Zr�#�o�!}�%3�B4D�pn\t���V͞؎i�sG0D��ڀK��/��r"�0�r%)��.D���u#�l<���`��MfNݲ�M-D�J���p���s�mX�1F�K7,D�PsC�Rj�����RLmXB%D�d�5mc�D��aiT�u:8}��#D�Da�H/6)bY�dݹV(Yxu�-D��Ԇۜ��e+���
Z�H�c+D��c[1N��A���5���R�j-D�xJ��S�u����@�b�``���,��h�4`Gf����B�f��C�Y�h �ȓ&4e�R�:�t�Bt���4!�ȓiW��
G��#�>L�s��)�z��ȓ3��Ց�B�	N)��ܞ.�4���o\\x��63X�p!Q��2����r��)9V	�4!(�E��
yI0��ȓN#�S ���(HG�ϭs�b�ȓM�@�y��/^��6"L�Q�ȓT��"��԰�h���֡�X��gX����H��O \�j��%g��ȓ.��0r��ݍ4�8�Q�<o]
@��I�L�Ӄ	"&^B���ǻ)�r���<�@,h"�L�\.t�%��6���+݆=s3��W���!DK҅��݄ȓ�z(��k���V��EU�j0���ȓ�R�Z��L�^��+��Q�k2(�g��~b��Y2���Mۉ\�����[��Ov�'	|�c)�*P�ӋA�1��Tr��,|]
g"O� t��v��,l��A�i�#�A�R_����)ҧ �`gc��Qq��a�.Jž�ȓT��1ٶKW Ĥ��@Ж3[^�%��z �'���W��-�:P�gK�.�p�'��Vhe����ȝ����9�bB�ɚC'B$XEi�3Q���R�( ����RO�tJ��BЅV�h�k�$G�n���BG(�<J��C;c��Ӳb[7L��09s*LO7/�I�QT�b�-��,r^ѳ'ɍ3?�*B�ɕ{�z�12LD�|��x9r�e�RC�I�f7�a��`� }�D�����B�I�5cZ����P9��S"S�84�"<�:��A�����Hy>���M�9#.�@�ȓC|��+t�/)<e@C��7hL�ȓ~��)��X9{���R��;'�<ф�J��,E�F)�prc��r���ȓ&e��[���88�£�8Mu�q�ȓ]o���1(�v�z���0rp���S��,�?W�Rqj��0)���ȓv�
�p��<@��x�t�������{Q����nU{��@�FF�����J���7 J%M��1)P ԂC�Fź]�� �5ݺ vNQ�a]�C�	(,�x�H �+��PC0!�)O�xC�I�$ޔreM�]J�s�OO�%�C�I��
��
�;.b��Q�����@B�	�Sh�H U��2d��vޟwu�C�ɐE������ ,B�2aA��j2xC䉏*hTŁw���x�ʴ�Z�}NC�	=<a��j�#9ZB [,W*�<C�I/odٚ&KиO��32j�>C��妰pb�S<(�6���'���e��&Pb���+ƾi�0ES���|m���Di6ʄD44$�[�oI0�^���>͌�*R���+�,�$%`��&v��Y�G�D���\�kڦĆȓ?8��(p�-^`<E�.��d��,��2B�ܻA������=��ȓq�*M30a B��r�
Ѭ��ȓ4ᐥ�$�G� ��u�s�x�\͇� xp� !�\��Ӆ�f����\6����?O����L��$�\�����I?e����$BXQc"O0�t��~�����L1}0��{�"Of�����x_y�3mυn(D���"O��ue� .��AQĂGT�c�"O�к%'��_�� (��N�;�>-)�"OT%���N=$��0f1=�Zغf"O�3�ɒ�}��%E��_��5"O ��g̓��V}X��ܖu|�1�v"O��h3�Ɨ$b(+����'U�)�"O���p��E�P0���s6�hA "O���1���!?@P��ͽ[���"OH�	c�$z���q��W�hXX� �"O�,�!FL��`@� ˭0@��"O���H��"�:�po��>:�""O&�h���Uc@��w/�uS�"O�9���N0�@V�r p�0�"O�K�b�g���9WE����	�"O��@��˜txs��u���:�"O*���e�j&ਣq�Ʌ:�xa�"O�X#`gE� & H�%�S���:�'�u�aL�ބ	������6D��2�gX�Fl�!�fG�5N��e)3D�� xk��+�:��Ç�'���d"Of%k�߃3s�l��On���"O�0;r��(A0E#�Í�5VΜ��"O��炍S��(� ��Er��J�"O�첗������*ݜA�Z-���'3��'���'b�'2�'�"�'=Ҹ���O�:�
9��pxF51��'V��'���'I2�'���'B�'X�)�w˗�c��] �Λ�c5��0B�'���'��'	��'���'}B�'���[���,8xT�,ݎjڌ�4�'R�'�B�'qb�'.r�':��'}��[ 
жO>^ԋ�6	��P#�'�2�'�B�'5R�'��'���'�0T��ˎ�uW��a�h]�0�4=���'���'���'b�',��'�"�'��\���l��Fj��JM��':2�'��'��'��'���'�]C@��'k�����^;P�����'9�'���'T��'H�'���'QlpZ�D���'���l1��'"�'�r�'+��'��'�b�'x�U�As}�IE���Z����'j�'ob�'��'k"�'�2�'d�ū� K;6\d�C�[�aNİ�e�'4��'���'!�' "�'D��':43׮�Q���jҋ�"dR����'�2�'�r�'jr�'���'Xr�'�8�[W�+&WV}c��C�H0��'���'-�'{��'���b�J���O4�I�;'� )��ܒW�L	geCy�'J�)�3?��i��M#Q$߼P�\�8T��4p+��۝'D�	�M�R��>��@$�m(E
,�$���Ŵa ���?�,Η�M��O�瓸�rI?��v��'O�L8��ޚdJ�v)�ڟ�'��>�3��	 ~��,�&�8.%�r��4��D�<����O0�6=�fQ���&mD�S%ʟ9�|�1fh�O��D|�pԧ�O��}@Ĳi��d��o����G[��H��D�<U��|��� �L�=�'�?��S�:��7䞘MA 
VHL�<)O4�O"��~z��C�8����Pol��d��m�<i�2N�>����?�'�I�h����!k�%��ѹ��ΦBx��?Aԡ
D�:l�|Bā�O8l"�n������G҉��Q���:(O˓�?E��'�Q15�QC-n0�f���*���'hd���D���?�;Hm�5��$&ZLɊ�o׷z���Γ�?a��:m�%
�n�j~�:�����F�4|I������G�ҙY��!&�|[�b>c�(���Xi,�򵆞>�2	�f+?�X��� �Ij��/ڹ��<�F�Kg�K�aL1SQ���Iڟ�$�b>�����v��*HQ�u�VNSϒ�`�ISy�i�/9H!��%UE�'8�I�{B�0�S�\�LQ��@Ż[�T�����	��i>��'����?��T�B�~Yʦ�  &px�BN��?��i��O=�'���'2�R�l𙔇݂t7H�c'9G� 6�i��	�!��0˵���U���+�ҵXC�?��XwBr������r܀����]'ۂ,{#�R���h�	���I����?��4��L(3�K-\S�1�٨H>��?�'QyA{�4����(S�	y��4��Iɋ���v��~ݞ��O�����D�OL���O���E"�p�␋G�-�f�20��\e��d�O�����������x�O�u���ʧ{U��e`
�a�h1��O�@�'���'jɧ�I�l3Hi��� �ֹ�"fS!c3Ơ�4#w��v�2�����jl?QO>h
�u�lE��CΤ�����F��?!��?	���?�|Z+O&�nZ���d��=Z�*��&.�\�.�	`y�mx��⟄��O*���'*f�I#Cɞ�r��	Ȫc�����O�;&t�t�ҠP�w��>�O<�T�sd˾@�$�5�ƄQ��d�'C��$��ڟ��I�H��k��fI�d4��*�%���0m_���?����?yK~��JV��w�����gӆ�a�B&4���"�'���|��H %�6>Ot�)�ݼd��͡��]�GoP�R:O�����?)�&5�Ľ<ͧ�?y&�^�2��Aϳ9^9������?���?!���dXp}r�'���':DݫSO��q����u'��	b%"��h}R�'��|�k�=-��b��GT��+�������9���K��wӞc>Q���Ov�D��:�:�#\?�
�#PÔ�p����O���O��?�'�?i�)׿l$P�(�>���+Sѣ�?YR���I؟Pk�4���y��V�\u���6I���1{�T9�yR�'���'0�d;q�i��ɪ}��<ޟ�l�  _�_�@���-="�j�F(�$�<���?A��?	��?��V�����b�$�M�ug<���B}�[����U�̟DˀI��r֦	���ū<T� ���:��D�O��9��I�_�8�ba$^�9_
�TBG3Y�Q"-@+a�Ɏf6��p�',��'��'�Ҍ�2lK�h�q��dϤtܼU��'�Z:���'��O��I����O�|b���+� ���i�^-����O&l�A�U�	˟��i޹��EFBF��SPqR�JrCRz��lla~b+�I��d����'ֿ� �%I��?���H"��8zBݙ�=O����O���O ��O �?ّ⨐�k��KQ���y����ܟ8�	��i�O�S4�M[J>	Q�̨<���h�ǘ"	���ȟ�䓒?��|:���M#�O@T!1j�3'\i�R	��wH)3��nd�9S�'1�'��	̟T��ܟp��M�L(�ç,,Kv�E@Ц,��9�IԟЗ'����?����?�,��٩���|��A�҄���)�'�<)���I��p��q�)*�jC5]��3U� '��9�k�"��TcF�-�M;eT�擶2T��)��rvq.���R<��(�}e�]����?)��?�S�'��T˦i�7eZ�L�J��s��"60|�9��`���I���۴��'����?��֕%ne�d���c�d�6�ͤ�?���#\���4��DG�{Y��O��	 ��ݱ4�N�;(:l��"�7uC��\y��'���'f��'�b^>�(R.�?u/���
���D ˂����O2���Ov��4�DX�����X�%ϧ?�J���E
B�8a���t&�b>��"Oצ��J7X���1ր��FAP�`�ʸ͓\|�A�C��O5@N>�+O����O�$H�6>m�qvN����<j���O����O2�d�<�F^�p��ȟ�	+1�pX ��%��7KÜ��?)wX�p�	�,&������q�ʃ�O�|��1�0�8?9�S�_���z�4q��O����?�`���2��t.�0:�*�c��?����?���?a����O�t�e�
2�;Ъ�8U��)	�#�O�8�'6�	�Mˊ�w\�m��o�o��h�e	��H�'��'Y�CZ0Mܛ���`� ��4&��ۂm ZM�0D�������J�$�)$�������'��'|"�'���r'�q	>��7�'�$}��Y���O����O��!�9O,��F��윁P@5����j�F}b�'��|����?>�MÀ��.� ��.�Dj@�Իi?�	� 0�1�OҒOʓ@TL����3���%ۥ9� <��?���?��|+O��'32��%X8�⡩�$_�bh�O֓¦a�8�T�O�$�O �$A�6��\���MP���`�I�T50]s +l�V�'�����K�n0�O~j�;^�=k@��4u������]����?���?	���?�����O�,�V,P��E�p��������'b�':��|:��q�f�|2AT�Y&lBA^���$��mU8&�'�����T=3�f��H� F�#��U*�CQ�N���A��6�3��'4�&������'0b�'P�M!WNU$�R��VhZ� =F���'��_�0�O����O���|2�)�/�%B4C�>���mY~K�>���?�J>�O�t�rJS*D�����u����JW '1
��"�i��i>� P�O��Ov]`�,����`qLչB�� ��O����O��$�O1�|�E)�o�	�VM�f�� `�ʭ�%- �y�^�P��4��'����?�`D�>�. #di� 9�L�U���?��_=B���4������]��ڙj�!��$�v�!p��T��y�X�������� �Iϟ8�O�D�Q�/%}>�3��N3U��{E�>���?�����?ac��y�*��xu�_�{���W
�F�2���.}�7Mu�$�AD���tYq��7i��;�cj���펔r��|��Uy"�'�beP"J-p�1��w�,H��@L)i��'�b�'5�I��D�Od���O�kt�ϾDĵun�-oBxt�c�-�I����O��$4���=\Y���Aѱ4w�sĄ�2'��	�c3�k@��eD�U'?�{0�'N�q�I+�T ���;[m�8�QHޞ������L�	����G�OC
':BE�L"w����/�Ba�>����?)W�i�O�NÜi�u; dR�O�6�y�-G :��d�Of�$�O��HR�fӜ�Ӻ���Š�J�&A�NH��WG�2���"�L  �O�˓�?����?����?��˘����n��$heM��R�DZ*O�=�'���'}B��ɍ;g�l��6��,�J�(w���'���'Pɧ�O�\5+0cB$�$4�QF�=1��	�FJ�z�º<��lD(<S���w��^y2�ƁD٥.��kP�`Yb�'�b�'��O�ɍ����Oޘ�sH߅ZFA��nG0\c��a��O�l�i��x�����'��(11�����a���&0KZ�X'�ɤ1����(i5`��;O�$�Er���)´A�	W05`7B�.0���c��y���ğ0�	�����֟���@�q.�H�7�}_�"�2�?	���?IV����ٴ������ˑ-��p���P���I>���?�'`XX�۴���?_����h�.|�	�b@�kcXQÖiC��~��|�Q���Iğt�	ß�*b7� h��-CzLŐt
�<��Zy��>a.Oh�D�|��LA�&.��!!=NL�q�W~b`�>���?)J>�OȌ٘��Řn�Y����Xܶ4�̘���-J�'��4��%{�KTv�O��vj��	��C�. 6���f��O����O���O1�j˓|���kA!q'R\
�jv�Xi�ФP��y2�'��wӖ⟜c�Or�Ė�&��ĉB⑏!�N�A���_Gl���Oze���r��Ӻ[@b��¤<� N�I�E��=�2ħ�2?/�I%4O^��?����?����?�����)LK~N�(�M'$]�$���1����'h�'b����'>�6=�\���/P�,�rOA��D+���O���(��i��r�6�i� ��Vg
|tزE��$3�� ��k�q�G�,\�C�J�IBy��'��өO fY�j>� v�TrVR�'�B�'��	����O��D�O�����M� �*�+ ��]ڦ�!�I=���O��$=�D�3]���(R�=��-��Kd��I�7N�Yz�AT$�Nc>ur��'�N��I&G�|k�E�=L��-݄j`��⟠�	̟ �Is�O�bf[�e �����!O*�(HN!ej!�>I��?���i�O��hZi�p�Òhcj�3�jXd���O<���O�<�P�nӞ��$�b�����q�<ߨ]��V�Y��&W�����4����OT���O@�D�,��̑R�ã!�k���_X�ʓ���ٟd�	ןt$?a�	�BŉW�i3!�)yW��٨O����O��O1�� hukU~X	�*��F`�嫂+"�|�����J#��WA�*�A�I@y"J_��I����{���5�n���'��'��O��ɛ����O�a�ą���i��T*Ŭ�y��O4�ow�������������1�W%����i�;3�,�B�o��m�\~���Q�t�Ӌ*#�O����m0�M�0k�[�Kò�y�'�r�'��'*���T	�RECU�O����S!i@���O���`}�O�Bf�֒Of)��,�j`J��
�).T�F��Oʓ5��ܴ��D��0�ڜbC*��=�w
�*��(L��?��@=��<Y��?����?i�?u���9E�X%S��m�e�Q��?�����~}��'���'��/Ia�ݙ�-F��;T풦���2���Οp��\�)׏P�&�di �@�#_�x�y��Ȩp��5��"l����dٟ(I��E�9��(��DB�ݡ3��1CWb�'�2�'<���Z����4^ ���O�(#�M���p�)ϓ�?��M���$W}��'*��"��R*.��m����J�j����'I�?r�6����<.��q�SJ���"�F��Ƨ�+!7���+#��IJy��'���'|��'��_>Ep�ᚖ��D�����Ϯd��)��D�OH�D�O4����ڦ���(��ĵ#�dA*�M3#�r���ӟ|'�b>�;�����y̓=q�����6	��Z�Kr��T̓|��;�`���'�����$�'8��ԯ����AYa�M�i����'���'�RU�TۨO����O��DW�Yi�)�"�="b$�D�dz�Ot��D}��'��|*��0}sp�_�,>�:������T�	j��c҉8IR��J����=I@�$W-�iAI�V��|٣B�w*X���O���O���>ڧ�?y%�R^8�К�ϹvH^}�GϺ�?	dP���'��6�1�i��0S�Z%1�:��&H�U@�T(z����ҟ ��-I��lZ|~�d����k�RM���;`�p����@��|�^��̟��	��	���1!���l�B V2�FXkՍKUy�ʬ>���?�����<��B�&����R�K�� �F��u8��Ɵ\��v�)� -ґW��ZK�Ӛ5_���M��	�'j��94.�D?�J>9/O.-�A#��y-����߰jj!����O�D�O���O�i�<��_�P�iUa3�C�B,6�YSD� )��R�'V6m%������O��$�O� (l\�W\�hs+9W�@� �K�:7m/?	�J8;���4���}�#��8B8c5'F4��1D�l�I����ȟ��	����:�fȁb�\���,�#85��B�������O�,ԧ�d�'j�7-(���4C��p�ǀǈ2�z�:U(��'�P��Pn�����'�����JX�z��̠W�
T�D)��eʠ ����z�'��Iǟ����ɞn��d�G�ӽ5V0���ƈ�
d���	����'oV���d�O��'K��`�&�BE'ܭ
CA_Y��'�l��?�����S�d_�k�� �&@�T9QdF?9t�]�&CڶDLR@:�_���h����|�	�+�u���%�-�"�%/T����Ɵ4�	��H�)��dy!g�j����eo�p�%
,O�N���5Ox�d�On�nH�	ܟt��O�����B\��k�"˄0��T���vL���O��8�`���Ӻ���I����<�ƊX+z�:Y��@�,b6Nd�Sm��<�/O��$�O
��O����ORʧw�ڰ��K3]l,���+F�p�Y���Işl��x�ş�����S�Κ�^�p6�1vN�����:�?9���Ş/���4�yBW�Vgzq[�@���K�d�R�'ez`p���՟KƘ|�T�4�	ß�[��w���0TaS����*լ������ß���ay� �>�-O��d�u��\����m�* ��L��l�t��O���O.�O��`DM�f���AT�E3J|�����ċ#�L�O�\��W�S�H�՟�1� D�p[t㉤Qh�u2�KD؟��	�p�I���D���'�x��%�#���a�������'mN듺?���r���4�*� �h 2Wb�k�"�h ���?OF�$�O��䙋h�65?A«�l�����c�? D0�E�Sb�L�"e�?0 �Ղ�c$�d�<ͧ�?9���?)��?�Q˚
��̢`�M$�zYH��А��v}��'|��'�O~�-�"k�F�Ч(�����K��p��?A�����Ir"@�d.��%rQ��@w�qq#B�Y��	L �q��'Pf]'���'�,��&�Rfv�ɗ�1j�]ʣ�'�'A���dT��	�Ob��ƙKv�I��3}��	J2�]	Nbj�$ܦ��?�V������ɪ,M؀*%�1(~�q㖠=ob� �MDɦ��'����E
�S�O�w��t:Թ�D:|�vr��B��yr�'Qb�'�2�'��)Lo��A�m>��d�eg������O����y}�O��%}Ӓ�O\YC�E�g5���c��{�nf�5�d�O��4�)3�d�,�Ӻ��%ڐI�xk��o�L<*v��,�����c1̒O�˓�?9���?!�J9��C��ri��@H�⩢��?�(OBq�'RR�'w"Y>�ٱΰ��%A"�I/Vd=�k3?��U�<�	��'��'0����^-G���y�H��1������'4a3v��R~�OZ*|��%��'y�E�a�C�lv���y�8k��'."�'F2���O�	�M�@i]�E� �o4� ��L�<A���?Q�i��O6��'T��Q5Xܸ;%��<d�°�s�S)�'��X�d�i^�I7�N�b�	U�x/,尶b�C���st��"l5�<����?���?a���?(����$]�}�|�{]��嗦$
�P�':��'�B����'�7=�\p "�9�훇�үt?�����O"�b>ͰB˦͓UuP��`m�G�L��4��O�j�̓
֚��i�O,�L>),O,�$�O@ ss�޹:gJQ*Wa�555~Y�"�O����O��<��]�,���t�I�}$����,kСK�d�GD��?y�S���	ܟ�'��+Ǖ ��)�o]v���%$?A4Dպ+�,e
�A�'#�&�D��?�U���b��1CV��8.�d��d�U��?���?����?���i�O�D���K%~� �጑�F���c�OЬ�'��'\ 6�-�D�O�F0X�*(a�N�Ig�i3En�.v���On���OjѰ +i�,�Ӻ�G�Y���K�~V��aL�U� �V*kv�O���?����?���?!�a{�c��I.?�a����13�Y�,O*�'eR�'GR��t�'��<s�aXY�
)�i�l	��!�>����?	H>�|�b��L ����Y�x��8��	/�
���4���W�0�~(3�'��';�	�+$���z�:A(�M�a������Iϟ��i>q�'6듥?�%	V`IF�wO���4�����0�?���i��O�%�'���'��G�gSؘ�� 2�`���ɺOd$%�id�I$�>�Y�Olq���Nҡ:B��9v�G�0?��
!�R(��D�O ���Ot�$�O���-��"0X��La�H\�2.�?Q���ß����4�������$��#�0�:��ês,^١3��|������i>%��W����'�d�C��\(�J�h�+q�$���,^uʕ�I�F�'v�i>�I̟����.!p	���[�2�x41�G��x�t=��ПD�'Ϟ�����O��'^A&�(UF�6g�a"	�6�ı�'����?�ʟ���gߚ\�.�@�,e�d�A�OgFV$�p�&���|��Ob�O>A5�A5n��XYҧ�&��|����?Q��?����?�|:+O25n�2�����ƶJ�hY���B"��IXy�Fw��DY�Op�d��V=��bhS�{A�qa c�П����*eo�z~"ꑱ��}�1,��5�p8D�$@
h��#�<q+O~�$�O����O����OZ�'UnXpEU.�v�R�7Wd幰V�`�'b��$�'V�6��l�:Р���L" ��#��'	"�|���o�8r�64O�1H���.fP��!��;%�<��;O.����?�S�,�D�<1+Ojh���!-O(\!�Բq� +a�'�r��?���?���@W�	���Q��p�o�'��'��듐?�������,���|�8,s�kL+3�DT�'��Yf��D2��w��d��ݟ����']f%E�PTj@aEj�.C���'�b�'�R�'a�>}�I�HDT��R��`�nM��ʓ�q ��I7���O���
�}�?�;�B�PulކkP����+s[@M��?����?)e�K'�M[�O0i��*��Z�"J�(�v�ۑ��Y�Bxz� ��m��OD��|����?I��?��i�ȹ��	ƀ��@�P)F�(F^m�,O8|�'U�	ܟ�$?Q����Q��L�-S�A5��s�O��>�)��6������_*ʉ@��D��Ѥ�Į(�䨕'�����ßD�3�|�W���#*�,N��D��lY����U�۟��	��I��}y�>a��|�h�%�	�k��,�u-��Q=��+��Es�&�D�X}��'#�	5L<�@ӒI3�&� ���D��Dґ��ᦽ�'W�
�MS�?q@R��$�w���J�#�%s|�X0���k�8Ź�'>"�'lr�'��'/�P}��A�$@@���I�L� 9tB�<a��?��i>9�I��M�K>b��%g��`"3-�P �q�!���?���|b��S��M��O�+p� Dh2��	q�.5��%ʳ,�F%��Ʀ�?A��2�Ħ<�'�?����?�ס�>}�����>10�B�J�?i����^}��' r�']��K[�< ��9H�:l�B�����n����� �?�O�>@)V��0��bBD�W���냙bbT�q���8.�i>�A�'�$�<�$lم&�h
T�A&�<ᒆ������쟔�	�b>�'�Z7�V=+ �تU�Y$\k�4zB�S��$�O���
�Y�?a�X�\�ɣX�"Ę�΅-rOrMr@㎵$���I͟�!5-��A�'7f�r!���?������#�Z�Bcz,k�o	�j��t1O���?9���?����?A�����	�7����áLh���E�H�'�'�b���'��6=�b�ڥ���l0��+��ݙ%�x��/�Ox��/��	јɬ6�{� � ��!�y��7blxpz��Y�v�"!�D�I[y2�'OR��6@�j����;yx@4�M��2B�'nr�'��I�����O���O2��p��\&NY��ļ
�^���2�������ON��%�D�|z�報ʛ;5��ʐO�|���7w^�Uq��\9�c>ay��'�M�Id�.��wɉ�#� E	��9F����Ο��������G�OM�FE�R�z5C��8b�Qf��$g�n�>���?���i��O�P�\ iBf�8kz�H��Y91���O���OV�K�,{�j�2���Fά?�)Ǎ��
[�͋*�

�Na�U�Z�	Jy��'���'gR�'$⎐"�����,
$^a�dH5O����ɿ����OF�$�O�����2t���RA{�I�I�Z�:��'�B�'ɧ�O騈R�&(�)���F^�p�7�͍#��v�<���˽8nf�IJ��]yBAE�?�~ԣ�ώ*tp��`,L%"�'�R�'��O��	����O���Do[�v(d�RWM_?i�\p�v��O�QoZM��k���Ο�������$�U.S��C���9/��]��"���4����=�Ra:����O�g�_�~pő���VJ��U�y�'�r�'0��'(2�	���,�.�+��
G��<5k����O���Wf}�Og�$i�z�O�X�r@ιV[�X��O���R�D*���O
�4���1V�t�v�-��p�ˢ[h�4�"PJ�̙r��
!���K��䓠�4�`���O����Rez�۶gX��]�a Ƶ���O2�$�<�^�t�����L�$P��mY�*A-<�ʘ@���y2�'���?���O�"��s���c����0`���zY��Z��	���BpW�`�S�&��_�&z^�i`�'L�V�<���Qxi���Iɟ��	ğ��)��Ky�Jy�hY[��ʆ	�l���C�!UΑ��<O����OT�l�x��	1�	ݟT���J5��:"�͇8�h|�`�Vş\�����m�D~Zw��*R�O�h\�'\P�Q��_�K~�͸"!�����'���ğ�I۟(��ӟ�Ih��K}[z���O��$��`�G�;����?���?qL~Γv	��wN4�iƅ����C��A�~;f;��'2�|���#]�NU�4Ofd���"
����NP�6=�4O�y��A��?Q�O3�D�<ͧ�?1�M�:�x���h!�A�7����?����?����D A}�'���'>f(*!-��iݲ�����	}T@s����N}"�'}��|BcX,���#�O3�L�zGnE��$�*N�����Њ�1�������j��O�6�^ �ІРDe�=����b�X���O����OD��%ڧ�?��䕪'P��Lî|�:��4L��?��Q�����$��4���y��� �q�1V@Z��4jD'�yR�'C��'�}���i&�Ɇ�,���O����O��W�mK��X���L��%}��Oy�O"�'��'��˩X�d�!V�2�� k��J��	��D�O�D�O~����J?�Q��l^> �v%ȳ� \�� �'S��'*ɧ�Oݢ��A�B%7Xn���أT[��kF�Tq,|J�O�����β�?��$+���<��bL9]�օ� ǽ4&�5�!g[�?)��?	���?�'��F}��'����`Ј_�*���i��~6d}C�'$"7�5�I���O,�m�('D��md��dEQ�2y�i����M��O��W��� c:������(iE�@�GJ}�f<+a4O����O����O��$�O��?IB�$�T��vN$A]����䟼�	����O���O�Moh�J�����f� �1�ܔV:8$� ����Sg�2}m�Y~����;�jY`��Г.�j�r�Q��$E�Ќ�ğ�r�|�\������������8E��B�̋v[L�X ����	yy��>���?!���	0K�B�j�jQ�'��c"�"��,��$�O��$%��?�3��W�o�Ds��6j)�1hVc_:#Л�Ɋ��M��O�Ɉ8N�QC��(.���"���I�h1�T"�lT���o�LP�A+D�Ne(F��j�X���k�$��DnV�TxA��+X�Wf퉴�J�o��5`�Yf��aW��-�dٱc��OH�Y2�y�X¥䆍bG�M �e�3m��ce�;�|�1��X���cM4LF0ѢK�Itp -9x�a(B�=?Wp�pf̀;Lhd�Ga�V�+���w��E���,n��ݻ@�R�,���І�Y��@�B�h޺@% �B�B�x=	�Z4_�E����-�-¶昄NrTX���g�4�1�i����$�Of�O���Ox�����Kr���po[Y��x�p��� �dפt���O^��O����3� � q�Q7F�x�)�F� 7��b�i!��'��|��'��,�3 QZc�98!'[�(�s�/ �L���n`���Iʟ �Ɇ��'H`��ǟ<8aO�76KL�KQ�(��\���H��M������?���4s�{B�BZRt��� �m�$�,�Mk��?Q@b]�<a�����O����O��be�BWiZ4�B%Q	/��Ԫ�j�f�	⟬�I)� ]�?�O�f� 2/�~L��F�Jv��k�4l�x̓�?����?����?���$�.V툍�4��L*H�@$$Dq�mZ�p��g<���?�O{M�شp,<I�U��'$�8�@D�␩m��|�ܴ�?1���?q��k���Hy�JR�����?I�K9�p��i8m���d�|�PB�<��U��R֯ޣ�H�����7OgFa!��i���'���'l�����O��I�]� 8�d�H&	7��@�*Q*.�c�,��OG˟���m���۟�	3 F�%�%�U�pn�xR�/z�q��4�?)�vL�IVyB�'�ɧ5֦
^n�9�ïrJ	��I���� �tyr���;2���O����O�O�<�w�̐*W�!9]�Qoߟ�M[�_�4�'���|��'�2f�\zb�O4L�2���Ԑ,��A�'��8�'yB�'Oҕ�dz>��Q/��Eb@�a��0g6�8�k��˓�?�I>��?��Ɂ"�~��t�����E�I&�a������u5O���O��d�P�SX�t�'�ҭ� �`(�� �͔�S�X\1VDe��!���O �� �w��ؓ�n-Zv��EN�e��bhnӂ�d�OT=�B3O �d t���'��5��ɢcRpP��\	�����F	������ON��/�9O�N' 9�Dkc���+���iU"]���˘%�yR�'�7��O~���O*��\p~�ߨm� ��mr�\�5,x	o�hy��'�b�1�i�|.���I�n �B� �3g�PDs�ǆ
%�Iܟ��	՟�Iן�������1�L�f��,��fi�4YN�E�'p��#��4��y���ܙ�a�v�pч3g�*F��6�M��?��?�.O�Sa���'f�S�"V/"ux�kJ�.@Dx"�}�����"?���?��@T�������8� ��__|o�蟐��XyB"�~*��j�)B�^�S��ٲ]�"�k��ǘ5�O�s kR0N������i>	��tغ��#�	
#z�����v��nWyr�'Y2��O�I?A�vM�%��*qJʍ�s�C�,t7�vJ�ɣґ�d�I՟��RyBџ�	�R#ֱ@�*4�æ�"\��ԷiC"�'?�O�ħ<)#hFϦ���)_��prf�*Cxͣ��0�y�'|�'S����OR�)_�*܁J�H?�� 
V�G(��6M�Oz�O@��|�����ʔ1�C� �õ�k7��O����8�\�,�O��'+Zc!�d�cN�tڕ��HƣD�x�K<!����\����]+�� �E�Q�g�J@�d�hp�7mȦA�$�O^�mȟ���$�ɑ��$�o<V,k��v������4T��]����ן�J|r/�.��p�i�6�i��K�@!jp��&&���O���O���O~�ī<�O~4�^aP(@5��?!?T� o�>y��W����!��y�'�q ) �c�Òj�*1ɑ�qӲ���O(���O�<&��'�~r�Y�� hh�)ԁo��L����M������?���<1��2۴�?��KP���G� �$���#؋	���'��n8�?��'�iY�m�dq��� ��Ӥ��5$��',��y��'���'����� ©� ���Kv�F�n��-nچ���?I��䓚��$�!��8�) n�BfP�!p�i
B���yr�'��'*�O�H�ӵ��0�#F�xT�%����ISv��?����䓰�4���d�~��t��@P�aZwM���� 1Op��O�v�Ӊ��i�O�t�!n�>Pr�Ui1ǜ��`�s�B�ɦ���vy�'�2�'��4��O��^�\y:6͂�j��A�T�m�<6m�O��*|��D�O&��O R�'���+#��L��.��.�)���?x����?���?�ǡN�<y���?i�nM�(L���Ϧ=I�Q�|�<Pr�:O��������ş4�	�8!�O�NΗa�mjeNAb��풁j3�&�'�b����y"�|X>�`�tӖ,9S�xX^\p��|�L1�ߤ%^�`k�v��O����O�a�'��ɗ0ȼ8�� !
�2�.��XǨ��޴o��Γ�?�+OX�'=9.��'�?Qp�E.(N�!7d�O]��@�j�DÛv�'���'H�>!/OR�d��$��=��1
���m6L����v�T��<A���<�voP�|
���?��b��PKJ���Ju���~#,PW�iB�'Q�����O�ʓ�?�1;%@��dV������d JM���'ڼY��'����u�'���'����yZwf8���Ӟk~�M`f��
�R�2�4m=��Fy"�'��Ɵ�����;��̏7����q�2b��Z@��7]����'d� �	���Iȟ�%?�ȝO�t�e�3O�ڌ���B'n��)�4��D�O˓�?q���?��'Ha}����E�x��4���h^Ċ�iԴk���I�P�	럴@Yw������Ok��q���R<f��,�%/�F�'��I�|�Iџ�S��(�s�򐚳BW�dJ()��L֩7Ʈ��idR�'bn4��'K�	�~R��?Y��1+� �R֩��Rd�B��]d��2�_�,������	�S�@y��'����na����� �:�$��2˛6��y��'�6��OV�D�O0�\R}ZwL����߹!X�� ���(�:ͨݴ�?1��8=̓�䓒򉙒Y���/�#N����dO�dK6iд��!�M��BZ���'b�'��'�>�(Olq
�
�V;��Qc�W����
��Ҧŀ�h���I^y�P>	��m>���	.N�1 ���c QA$�_ e�2��4�?����?	�3��Wy�'/���Y�0#���3]��͚D�" ��ayb.W�y����4�'�r�'�~Q�K]�{�V&O�]�*IS�(�b�d�O:��'��ޟ8�'�Zc�d�"���	3n]b��Đv|`m�OD���<OxI�D�O>���O@�D���f�����iM��{�� 6G�0h��i/�ꓓ��Ox��?y���?I��R�.��$"�Ex�X�En�(���5݌�ϓ�?!���?�L~�5ܟ<9��Y�?�Va�垦d]T�L<������?����c��#,J��!�p��+�T�8�#��<1���?���\ÉO}|��2�4T��ٯw�|ڣ�����@��i �|��'!��S�yҐ>q�M�k*�򠃔G��M�Un�Ŧ5�Iԟ�k'`��	 ��I�O����O�Tʄ��9�ZyB��I�8.�#TŒC��ӟX��){�X���j��e*�\?".2�h��I����#�Nʦm�{�8����MC��?���?ф��<�V��l���B�O�y4����h�(�D�O�E�9O��O�]0X6M\�C�б!&��`s@��Ϳ�&�'`b6��Of���O���L�A�ީ���]�S��(be�$,�-�i�h|�c�'��';�Ӕ$�����dh�O݋Bw�Wϒ]<�$��bM�M+���?y���?�5�x��'���O�t%�z9�����,-?ֵ��iD�'�R��'�^�8�'�'�2
64��k���<f&�S����7M�O���D��ǟ���c�i�� �#Ί-���zCZ�k:��tk�>�Я=�?�'nA�<���?i����=���`�K��e(Ύ���7Mu����p��Z���t�I:-b�0�݊��"V"ݷg�Th�t����T�w�d���4���9�2MP@/�.|&�0�7�֝y攤)vS���I䟈'���	������<�'S�:�C��GD.�@[a��A���<����?��f+�O�(�'�?���ȕ�܀�#莽;�rY�+	:v&���'m�'���'�*R�'-�Z�2@�,�"�9�"RaT�9l�����I�������������Ov���*X<��Dl33s1j�c�H�%������Rсg�$$����C|0�i�8F@ա*�/x�BMm�y����韜��4�?	���?9��o���6"��q��*Ir`��e(�v6M�O���ֆ4����9��|�A�����B՟h�f5QAa��!��(Mg�2������@�I֟��M<�'�X8Bң��\Ƥ�+�C�|���h1S���	m��|��M��<��2=Z�"#���,�Ā#DA^`�H�xe�i{�'��'W*ꓬ�$�O��	�>㦄X�� '���@�"�(n��7��O^˓q|f����Qͧ�?A��?7��?p� X�3�,f�ڱC��M�1ڛ�'BC�>A+O���<I��CU�ϰx;�K�d/(iF=���K}�)�y����r�'"�'����u��z����'�ΫD�>�p0����MCf_���'�]���	̟����B�81*C��9�S@I! ��q��w�ʃD����I̟L�I�?=�O�2�S�jn�̠a閩8ڔS�'��^?�6ͬ<������O.��O���;O�x6��>Z�R-�V�W�(�|��P����O(�$�O�h%>]�����>f�4��SG�NlH����M�¤n�ޟ��'��'z��V��y[>7��ǖ���n�9Rf"x"��d9�&�'��%���y�'ƈ�'�?��?�qLJ�Y�ޑ��@���m[VL�+�I柰���p25!a�t��yB՟�y���|����0+E�r�dH#��i#�,:�')bw���d�O���&���>��4�@�5iwUD�r��8<�0n�՟��	�T��������OB�'Ds,5�;	��`���f�*�Z�	�:΂@nܟ`�I��L�Iҟ@��@'?���H�y�D����^�.l(��G8��� Hh���!������g$/+��b5؇vjԠ�ҁ�M����?����?��x��'4��OpL��[9�sGbģ6"�H���'r#|������Iӟ���̚�v�$�eE!?ke*�7�MK���?�ӗx��'�|Zc�r0g,ƴ,i��B��҉h�r�}�ͅ�y��'���'&�c�� �m0�b�% D�wOn�n��ē�?������?��&p0�F�U�?�ܱ��F̲z����-�<4$��<A��?1���'~���)c��j��A\4��£�+;)�	ڟ���S�Iڟ��	"%+h�h�:00b��_?,�1%-�D��t{2OJ��Op���Ⱥ�(�(�'�?���_�y�,(
H.M�8�bS�$���'U�'H�Y����:���ZZ��S*G�|2%kWa�w����'.r ��y�']*�'�?I���?)ea��o���e�W�r(������fQ���'^�)�ɟ���?7��=NC�y �B��~ �ѭŢa��&�W�pEB�'"�'gb�'Q�����͆;^) ��$$]�SN0�M������"��ӏ=""7Mǰ��X�PΙ,��ZAǭ��V�'��7m�O���OJ�DEy�̟�� y�a&��CԶ�P�a)X� dҷiXl	
��?U
Gek��	3�¤��e�Pr��;��o+��:�4�?	��?��!d�O��$����QB^�d,#vD�j@(�b�5�I*Rl扶2��������؟�Є�I1|��|�7�G�mӒ��q�۳�M3���?���xB�'��|Zc1r�iV-�L�x08�)��9:�{�Or�p�2O�i3&6ON�$�O���%�tc�3��=rF�ST�"	r�)��MT�d�O"�O�D�O�L�J��_4&h[��"��x�#�	q��]	z����O����O$�ɤ|z�O���ǒ#v���S
D t�HIش�?Y���?�K>Q���=%��F$� Ċ�c�09T`t��IE�K���㟔�	ҟl@K|RW?i�	��0����:8����= ۴�?����$�<�tO��O��@K��<nm����R�*��i3��'f
��&�'��Q>��I̟���Z���RD��3����w.+���ē�?9*O��ّ�i��WǑ�;*Ѡ2��?�� �"�z��|)����#4Q[N�g4�x �
ʜt`I����+Ԭ�؇!�f����уN>%����7H�!35"���޶&I 4�ьW�O��I���+%+�=�R�E(	��Z�J�+'r`�s�ٸ:qp c�C �<)�ER F���N	��|Ѳ�JjL��u��1�����'ߨ1JdGW
R3�|p K+�DDzFɍ�m)lAy7χ�o��r�Y�m����W@�m�h'M�7���ʊ�q�9�͂�{�l	�H7@�Z��E�E?�s'��C�R�΂(kF�)�!����4�?���?�,Or�d�O20��ꜧ����GHԝW��	q��ʟ8���F�L��Ex�,ƈ&n��	�m�|h�e�S�%\d�wf޹5� ���s��Q#!C�!CGv	R+�?�=�rj'%ҽ�4"˟]D�ja�N?1��U�$�	G�'��BR�J��?%h6�#��:�B�I�� ��9,���S�
jP�K���?�'F�xC�rӸ\�D��
tUZ�P�hP�i������O��$�O&˓�?I�����W� ��/H�$Y�֪Y$T����+�%	���g��/Z��y��͸=�$���۽{� �qS��`a���ʫ$$��g �xx�����O@�Dō6�,)�D�[N:�:�gZ�*�6�=����V��T�*UH�"0 �!��V�!���ك�׬bvLi7cW�\��$AB}2R�XCe�����O˧˚�x�	p�|���h��h��?����?�ph�,*�F��\�H���S�d[�X�*dM�+���#�A��(O�H����K��|Bv� f�'%�C���ac�]����C���Fyª��?����Ox�1��s̐�+/D�L���X�'O���U������!�6�DL�:�0>YC�x��W,k4���%�KG x	�`���y�&�aӼ듕?�L~����?��� �����՚�#�� �y����0��&,2���b��S����'�"��IΙ۴U�ecAZ0h�0���&�1kڌqԧ���ن"X�˄ˑ���	K�F�(>�a(��'�"�����O؁�2G,��Ĩ� E�z�J3"Of�r���B�IГ@�%��l���*�HO�S�|%�L�F�N�o������J����Pr%�!�Ms��?�����O`�D@7O���0��Z���Bm^���E���}��\V5�T��o�[L���~�N\���>���l�pFS8��9�)Dv?�%������	�Z2T�@�C$:n��R$/
jrC�	!^ Pb�#�����G�n^V����]0�I޴(1\<�3$ ���͠ ��vYZ�����?����d�O���k>A�$�O���%VP��ԬӔQF�تD�ƪQ��|O���d��[́�R
(��IV��|��'�?y��q�0a[�ΝA�<-f��&{�L0�ȓ Ѕ�̔":*�]�� EbD�\�ȓ_�:�� ޤ�{_��(�F��<Y����&�Rxm������|�� ��(`fD�un
�$�yR�'KB�'Y�8�'�*�O�S�)rL�ؖ�T�䁢@%O�Q�l�<��+ۡR�Da���w��t0��JsII`�Fz�Q��gH�O0�$�O�Ĩ|:d˂���h�N�I,�MA��5�?	���9O�P�Ģ˜<{�}���X(��'H�O`Xu��
_U� ��B֥; 2�
a9O�� DM���	ݟ�'?��	ڟ@��%9��asD@%��{tKS�fp������ �<��O����=8~�8ye�ċ*n��q�J�Y�#<E���E\��J� ΉuJ��֫�I2�X��ί�?i�y���'���1e�,�����̆w��Q��'H��&I�<_ꨁ4�E�m�x��������	�S]V 1I׼Pr��l�|�����O��C����i��џ,��Sy��y�C�W���Jk,@z��k%�Ġ�~!Y!��>� �y�T����`a�:{�pLj��OnÄ�'��	�Ȱ+�
���#X�D��!I�'C�]�����=Y�p@����@ F&:d�@)��<�d�3E� =#���=p�Q��ϑ<3Y��"|:��ļM'�����o�=yB��o��pR�O��E��'��^����4Χ�a�I��xAVʕ q�ʩ��^�;�2!3dO5�O`��Z�����F(}x@u���[�0Ų�a6�O����',rv]���@�e��%�����yrm\

��Y�0���VYB|�aD���y�o�
d�\16EȊJ�6�z S��y��5�	��dz�4�?!���#	BP=�' U*ixdS���m��d�OD���O�ԢU)�ODc�ʧ#��l���	w:4��`��Q��<Dy�(����Dݡ@J�*dQ@9hG���x�y�c�I8L�D ڧ	�Ą�%nR�Y��
���5�\���@�#	�`:&H��ΊLu��	��ē�pJ�$ޢk���D��z��$ϓ>�j���?I��䧈?����?92�U�wF q�)���Hɺ��C�+���i��瘧��	[d�B�$��H���P��s�n����2�ͯ*�ְR��οl�j��d,��C�����'Jb�'�R��O<`�ŏ�J�>���ţ��<x"2O��d!�O���U�a�lAѴ�=y�0�B����HO�i�O��C��3��@���q���BR��O^�DN�b�=o���@������'���'mA�W�0n�B�cMS	���q�'#V��W-�;_�a{"˪�n�FM	'��L�����~B��/#
0(��'�  ���*��+D�>o�M��'
����'$����,On�Ĳ<)`"�>��k�ʰ�씘���s�<ɒ��3,�$L	�넫+k�m�P�S����'��/Yb� l�;$�b�Q%l�.��!����;����֟�	FyB�'QB2�$���'���+m�
Xh�I��h����@S/�p>)��[y��C9Ko��c����.=0��p>����8�I�ᐬYG��/8l��N"N�fB䉇	��D�Ѧ��=�0�F � h^B�I?B��2 ��o6�M W�����	���'j�ER��
��O(ʧ`>� ��*�<ī0ɦ=�l�̓�?����?Y�/˒�?��y*�T�!E\v¹���S�R���+���.��*t�YV�0�����j��D:f-�X�'�J�	���h�>!�%�'Z���1��&ib@� �"Od�x�.�:
3���e�*`��L8��'��O�da1`��RU1���>p�8u 5O���Bզ�����$?��I䟸�	 %�4�cU�B��Xa��+,~LAJ H]����<��O��cx�bX�S���f���*L�	�"<E��M\�$���3LB�!�W0\����N��?a����O>����� CVLO�A*dQ��[g��$�O������G��	2��$,)i��϶W�"���?U��ˁr ��ÖS�ACJ�򥉝؟��Iu!t��4�?I��?�*ON�d�OT ��M7Ӑ�ѡ�@�g�t8���O4����'��J��Mz6�C	�Q�՚�'(���a��(�NH�3�-�5�H�P�0Y�vFr��	o��̰ӫ݇&�@hCm��U%<���1D�0vg�A!8�{�-�4]���獐��HO?�	�L�좠I_�Jj�5��*;��B䉼\G�p�OؓJyF�1��:6\lC�I���Cn��j2HA�ET&M`C�I�2�ƀ����W�(!J�l�Q�LC�I��V}�'*ʹ9�R��wHM��,C��02���O��X�p�3DM'8�`C�	�v����4�إ�0�QP(';�VC�		 �`d	�".Ӄ��O+�B�	C�����;b�┓S��rB�	�c�f�����nZd��5��2B��B��&^F�kE-#8�[�#I(j� B���`��5�ŵ%���h� R�L� B�3yxԁB�!FБ�DR�g��B䉬0g�� ���)Q�A�ae�f�C�)� ޭpb臕'�j�*��	��j�"O8���d�S�R@�F� xH�Q"O�4�u�Z�2�,�[ O�[%�5"�"O��
��ů$)��p��G�m �c�"O&����I-f�
��������"�"Oj��.�H���"��^%(n<u�"O8��� �3@�P�9x]~�C�*O:��V��>k։���� K�)�	�'�<��F%�l�,��tn��~�	�'�
��&B�r��C��>�j�;	�'�M(�g�>#0��a&�\�0	�D;	�'%��H`�ͧLL�2�Y;�D���'�h��a�nzQb��-�����'�P	�ѯR�&��.U*����';\\s�,ڹ1��!����=(�Lj�'j�h����6Q�h�B��/ ���
�'�ޱ0C�a���"@ �G]�*
�'������^�h���ųA��]y	�'<��Ê6�`$s��A�f�8	�'	2�k�-Gyl��H��;�d�"	�'G a���NG��E��C����'^��x�H�y��W�ȇ)���x�'x&�i�)�9W����S�!4�4��'���X�oE�9� pZ%!O�l7$�X�'D�ђ��=U��D�_���)�'� DY��^��qY��ҎL��4��'���JS�˴[���*w��2H),T�	�'C塜	W�ش�&�	�0h����'�-;ң�((@��8�F_9Q�Bx	�'q�CgB�j�"��5k�8�6�'m���Vp��I)�>Ӽ�	�'D�(A�n��q���h�n��	�'D�tk ��"���T���v=��r
�'F�Z�a͙�6u�TD�p����'Sv�í��0����3`�7kp�D@�'��T��-c���I�U�f�\		�'&@�`P����,9�NBh�,*�'���󠄤HVr��Cb�����'�(���՟U%��7cXY���'j:��!H�8"�آ7�Q�Dz�C�'5��p�$�!w��%�����ߓb ��OB��
E�Z���gH�1�NPk�"O&ER����?H����[�e���J��X�����X,2��0c2��i����"O����όQ���Z�Ô�4�c�ݭL��O��}�sPҨ��F�	`6E��(!r�:���x,�C#� *�d�a��M�B��I30:�!����H!�5W��+: Q�
�S](���Q���Z����P�Ȳa!T|�Ѩ� ���ȓ�h4�R
�	^r���XN�pU�?�B���~R�)򱟪{�F� ����ь1D0��V"O��ۆ�ȍi��L"4IV�d
��H�i �D�d�����DZ.P�4X	E�� y��I���D�!�ٌk[������.W��j�U��1O�h�E��p<5���K6�����+B�M`��b<1�����2Q%��bq��uf?Wn�X��&,�X���($�~��NAԍ��/'OF �c����'�\��AkgK&��Iμoi��'�>�3���]Vɉ���%i$���O���A����v�2��
!�䙕����"O.� 1 H�zL���O�,E5�<�g�D���Ћ����r���)\ۨ�����y�&��*[&% !���	[�@���DTL���;Q>b�Z����'��=���I�(����\;N�tB�c?}AR�<�,E�B�(����L={��u@�k��� �4��KJir%�O�	s���J�N^�|7�e��.G�/q��2�f�Tn�4D~�隀p��(�~�PK��H�>�z��2L@��c	�t}�5��Sn.:��q�'�6`�������Ġl�'l�*�g{*8X�����oɄq��d�V�2(f��4��ܟLc�]��� ��v~ʟ�@3%p�%r��%�
�d/)>��l9�OH�D,� K�zS�:e%�0����ʅ�rbIsg�'?ʄ�v�'爡QR�P/S����O�
����\�ϒ% �$�r׊�T�\8�=iAM
1��4b��'=, � ��[�I5��d*U.[�jY�Yp�V2�R�dY�e�����Q�Elt#�#U?wQ�<v���9E�\P�N�-�Y��%ؓ!W�H�W��%5��v�ex����_�,����-!w��sN� м��A�'�F��Ƨ�����ef��q.:���1�:���dĺ/�x�;�h�:�6p����0tDy�
�=�8�B��V8z"<x����!Tx�Эܔ�R7���KQ�uG{�$D"u)3���x ��(b�B4�~bS#�8P�B��
��PRf]'��'���[Ӂ�)0m�D��*%*i�N<I��H�!�Y8a�R��:&����v銥S&θr$M��#�XI��8�]*�@1��c��T:����Z(ӡ�43�(!8��_�ɚ��ɍy�`%�#s�60���B�-��ܚ�FP��~���88jP`���35)T7��>11!D1�n�����3�tiP�L��yߔ��P�N:�0=Q�Fܜ/JJP*w/��]t���J1 �t�j�dޛT΄u� ̖b�'
��PEP]2$��.�!2��'mD�R��0_�`�3�� �BС�y��"B!Bѣ�ND�iX�1��'�� �Ƅ��2�AB�T 6_^<S��)̨)Z$��0d�H`���e*�D}2�^N���V�c��u��d,��$�	ߡ�j�8�O�?��y�q�\0��gפV.�T�G!7�pL�S���Kt�ڹt���F/�j`���o[_X��Q��ϖ~	NP��ѲFƾ��g�C������x��̱�)� ���Gg�`�����Ћ3��<�&ǜ
>�dbm8ړ!��:��\�uO��3����zY�Y��J#���r%D&V��ybNI5a�(�$��{fFY!(��
�/n�BePeM.?�Ua2[Y~�0�,|�SG��.'�L����A�����O�5���pfĄ��~�G}R����lY��4+MV�rnQ�<I�&شq �M��lEY~�)M�m����b矪JG�y�g	2*�D!�����k����p�'Yq�W ��9��Q�eLˇgFuȓ� ��?����O:��)�5���� ք�#!��4+�PZq$=�Ox�[u�èga����ukf��U��ZYj��`%�Tp�'4��J%��O�ၤfݬW7
����b�K�'�E(;_�Ѹ�̙w��yӎ�$/R�<��
(L��M�u+��so������˚�����ʁ(�S��'8�hT(�;z+���G�%Ȉ���䗍,/��JP�J)�leeg��	^~�����D����&�F�&X���������xժD�c�m��j_�|��#��-J�:
�Ӽ�Q�� )"%X`��`�\d�R���<�&��OhJ>%>��ƭ������N�G\:�qL�F���yv��2��B���9���0��x��C�QG$�c���'�-Q��~���r���?r�LؒtnҊPiJqP�A_
���̄U!���/ �Ji{T���RJ�!�ō��B��B������h(��
T8j���@�Jh��|��ɠ���%�%lՆ\A���
)�R� ��x�I\yר�΋6n�J�	�"��0�����VQl��.��<9cM��ą�'�L��'Kh�����l�~�(��'x�����h�n�*���4J��p�E�%ډ�#�ߏJ���.��Yp�'b��@��$Pq����U�>��L��z�ܑ{ዕ���IE�v���-	��4mLdh����W>X�8�b̰i���28T$�0��o�q%�#:���*�K5?! �Z���ϻ+J0#�!V�|Kv�+��k1�b�bD���ٙ$_P �F�ߛR�J��?}C�X��ٖG! �FՠR�V�
�N,)���zH<Ѷ�Z.^�͹uB75��"S
S�Ġѩ̾o�I�x��}�'��h�����~�V=K��X�7 0;8hh�ĭ�9�"��2?0xH�D��y9"ԱXƲ���H��aGJ<#�C�PFh��Q�$Vc4��*��Ė��9V�	���'D<��ƋG��P�x��W�O���A�y�V�K���B��+<x�8�U�W)z��`@Y:�yraKQ�4�c" �$Ch�a픁���QCf�`I0���!\V�y&�9���f��>ᬤ�m��~�d�}�
c-Š,C���œ<�hO61��+�\�P�4.#i��M��c#4��r�)C��:�� iZx��	w; �0����<���5���J��K6h/�J�2a��ࣇ�( ��Գ�T!�Z�r�eK�(�J��@cd֗F��A��[������ K:��QX@
0�'���7HB�+��I�0�"lXi�Ó��\�D�A�`1�BK�F����1q0V���@�|��&m�)*N�k�?[Pu�c���<����m�0H��T+u�a�5�b~r����ôc��@�R��&	�I[�DY[�l�1qJ��H��Hb�@��&{!�� �0�E�։O��Y	7�F*H�2� M!]|z������03n�Şd�'̒�c��/8��t2@�I�{E�y�'y�a��C&�pU˰����8v��<!�	V�s�ڵ��!�<���Ak���6��$m�m�#�C�az�2O���g�c?� �l����h�/�fb6�l�<Ѳ��'V�QYgA]&�l�QZS�'ɰ�2��L�O�QSo�%F.�yU-A�E}<�
�'�V�KTb8S|�#�D���R�l��@-v�s�'8�g�B�g�I&l �����-殨�A	N0 �BB�	4j�ap�D�?z��VQ�}d"��7�c@��!'K��p>y'!́�^;��\<*�j��e�j�ڻ|\��$��:���O�6--?���
tI5C
�.(�����N�!�DS�ސ� �9L� m!�aǉg��w��!��̟Hju��4�U�/��ϧ7�X,p"���>��yR˄(JB���~$��ɏ��`qr�
�4���ߏ�M0��X���M�d��L<!W�B. 伳��V%0ޜۖ��Q8���s��_1OR7�F�`�L�����A�%CQ� D�H���-.�VтG�ٱ����dm �	�g���>�~�T��4g�`���2�n� ��@�<�0��A��@�U��0z�����Od�<�a��	6Tqx0,\)z�4(b�__�<�FjK�r)��8 aJ"N�0�сWZ�<�����S�$�R���0��E�7Cq�<�G^<D"�TLE�G�Y�D�V�<�&�I�!��t�!��?ipUB�#�O�<)�Ŋ>�8�H1&�)�.��U�e�<���I�N4��#sCf,���h�`�<��e�����M��P�I���C�<QA�.xɄ��b���"�R�d�<a7���:��YV~�eY��f�<���rg�p�uդ'�4�hb��y�<ApQQ�I��k��6�p�<9�I��QRt�#��I�؈�D+�o�<���u��hT��#M�P	��q�<y�ƨ]�}���Qs�#�w�<���q�R-b�%S�|��lw��^�<�a�4^�h�@4ٱM�-U�T�<9Ԃ�/��MS�bP�Un�DA�J�<1��4,��5C��J�x����M�<� MD�S��M˒�9X��9�'�CF�< �ĕ
zΝP"��z�漀׋�i�<�VJK;:�(p�E��;�����L�@�<QD�X�'4��A2L�Q���3�&GS�<��ĉ>p5
7`>6��9㥆w�<���Ht���8�*1��ؤ�i�<�X�z]F4qaHӫ�6���JRl�<Q�/M���(`��i���[_�<�5�6�>��b�{�J��"o�a�<Ԯ/��Q���o;b4�\�<)dF�l�X��e�l�����[�<s�L�oN�]Q%�C+,�*��_�<ySn�q�\���[&��$�[�<i��/�PK�!Kl����K�<�l��RJBq$ȀIGj��I�C�<a� �l��B�"��A���1�k�<�G��1���Bw�i)t\�bʅe�<��-�t�10HLN�ޜ$�F[�<QS�.lͺP��l�a�|S�}�<�eK�+؈�h�l�m��IP�k�@�<Tb�,}�$j�B�/>����oGs�<�� �0��[0e�!� $�g�<�6��<J8�ki�YX����d�<Q���DK晠`J�(r8��V��i�<Ya��c5pՈ aЏj	֙���e�<� �!�F���\�����C�"O��"��Pc4c�+*m |�P�"O��c����,~��%��u`�3"O���pB�|���Qt��%� �pe"O�TQ§Ɯ\Jn�;���-�^��"O�u)A�9g����9`g���"O���T��7 �Lm���T�>�ƥ�"Ov��@dْ)�(uKf,E�<��;�"O��d�T�Z��P9F+D�"w���"OHq�&��}���J��Dmha�"Ol���O��!0������rh�M��"O�`���U'�4 �ȝ*V���"Ox�W��%�lq�6ʜJ?��;�"Oz��]%T��z&	��2��{r"Ol�V��?
�4�#�_��f�2"O.� '�)1 $��F�<[ŃU"O�D���l�)C�4k�9�H	��y�)nD��۷���2J=�T�ʠ�y�G�"K��P��N
~	$��S�y�R	pd�p���G�}E�$c�-�y�*_i��@zwgɇD�`i#�/�y�$T�M�UY!�;AB(p2��/�y�ϑjT Ӫ��,�`���yBH�7�NԢ���T��!H�yrmU�pkRҔ�P���$D�9�yBg�0xIP��Ղ�w���B�?�y�m��?ȍ�n� ^�5"$L#�y�+�H��Q���{:�8�v����y�I[b�֪	#s����A	�y"$�`�L��7(��d��|��K]�y�R�Y,����C H��腕�yB臕/jȝXGHB���(��я�yR҂@�9�)�w�����Α�y(Y�z^��P�_>o�*lA��E��yRI�MKzy`'eߢa���
熇��y�[�o.�BRN��t	5J� �y��<�\�y�!
� � @@D'�<�y"�Ԯ~��Q�T�P�~��q��i4�yr�[�&c8ua�-�5u�DX�W-�yr�����r������@]��y"��8%��x�M	h�hbE@��y�!Ww� h,U��÷���yB���P����gg��|����ح�y�Fߧeʕ#��� _�:���^��yBE�A�Ή[�BΜC�Ju
�g��y�(�;&c�q�hA�4�
*h6,{�'ׂp���M�$�"L��Kl��h�"O}�۟r;�����ʠk!\12�"O�-�L
�� D
�U��as"O�(�Q��*V$C����Y3����"OX��e�6��P �N�Ȕ��"O�m�K�"��e���M�W�1�r"O�I��L��7Ϧ�;�@��~}�	"O��;�i�,ꜘX���:DȾ\�"O�ݙgΞB�y��\�:R�;W"O�8��
}�dY���i��h�"O�h�à>ӠÇ��3�z��"O�M�ƌ]*EO����#���Ҧ"O��WBS�}��T!	>��@"O8�$�"h��X����"����"O�I��p���Ud�<CO��3�"O�1��L){�H��`�ѷI�*�ڦ"OL���"��=��Jʻ��� �"On�	���Y��)�a�ײ&�|�#"O� �]
o��a$��r�̤Z}h�[Q"O�a�EJ1u����̽f�����"O�%0+��]�F`�j(�z�"OX-ru�/)��ST�X�NĦ�k�"O� �S4RZ%Wd~�~M�"O�S��V;(�v`��e����d2�S�|�C�F7��e�AL��XǂB䉧��pa���0}�� ��eV�aobB䉵t����R�C<�� ��;�B�	�M�����Ņ]%�<��aE�x����>٦哗P�X,�e�?�`%@b��p=���ט^�����菔��)X���b�<y�#L;Xbfb%�:紬�B.�^�<9���(\�+�"|JDKs�c�<9�*����]��!u,�R�(�X�<a�b$}�Y���H6*TI�`��P�<��cȎh5N�C#з[4�( � Q�<�"�{i����eܜ-�r ���.T�P���(�80q�K�0)����`3D��)�E4-�85�7��C�����H.D�,��!_F�XPK�4����.,D��!���)n��0�w�N�l܂���>D����N�g 2t��-�;+\T�sP�:D�,���G'�`9
��B��U���yRo)5�0�!�fR�}�XI�,��y2$��n}ȓ�8sM��z���y�D��4�y6e�g
����h<�yro¾t� Dz0
E�W�zȺ2-��yRǇ2(�t=Ѱ�@��In̰S�!�䃽4�tT��m�Fzq"	E!�X� <�����C1uP
삦�ݘ!��P�%^�I#Iٸ_C~�p��ܞ�!򤕔��Vk��r1&���̳w�!��9�1weWl%(K�m��S�!�D�=f��,9%�{����Ս�8u|��/�O�z�lA������I@��:Q"O�l�#Ɇ'*	9�Bk��%���"O0܁2�O}c���i� \k�@�"O�$�I�4c^�c��!s�A��"O����ΣBQ���6S�UƐA�"O��U��^�,e����):O��`c"O�� �H�jf~���BՌJ��	�"Oґ��P���!��k�����C"ON��cA�L�a�ȁ�0�5�"O2��P'R/V��{���&"��t"O1�%�R�.V��)�G�w䰋��	\����Z�:��Xȱ��3}:Re醯Kq�!�$��@<BP/ǣ|��p�O�m!򤝇O�x�8b�f�A����7Ac!�ė�W���I�Rc�r���G=!�D�J +�gŌ!!���%a������Q̓�d1開��T���s� �zA͇ȓB@&�`��<`� h�� #M�4��ȓB�!��
;���s&B��>��ȓLj�@���Q�<AQC�ZH⠆ȓ����/�iDb��r��C$���38[��<j�ldP�GF�x5��}T|�#�M�:F-���тWڴt��IA~"	��c�ψD
ƍQ�ޏAu�C�4q����	+c��4jU��	!�C�	��~�9r���p���(Q����C�InD��$�E�4Y�x��GR�;i�b���'��~'$�{n��gǙ.�*x��Ga�<�M%&�t)�ؽM��hk�e]�<� �t��BY��(7��.f�l4��"OzU�q�6�vyI�i6P�4"O@ܱ�.�be�#ٲ��"O�D�g�N�9Y�h�w�C�&5Խ��"O����()x�2�i� w<�T��"O�E�0ɕ .��鸕�Ҭ3 ���"O
4�U�R8U�(�s�&l�4Z�"O0 �+̬Ao��ӁU�Z�;"O�hW�P'�|#��$U�։*r"O�j��� x�@,�E��6�n��"O���҃R2��9�MLJ�v ��"O"�!UۗW,C�k�Akȥ��"O����ݔH�"1'�Ϟ1�X�$"OZ����._�&�����7\~x�i�"Oe	0�ȑ�������5�-:��x���[���OX������2�'��A%�4��'X
�r!���i�*m��K2</Hd��҇�HX��b� �06���	� �!7��e���0D������eCQ���qw�ih<ib-A�':�2b�=5|����\�<�A�W٠�l�lF��Q�X�<I���r�(�"�%H�?�����Mi�<����w\���O��H�c�96�!���hV�`��i0,M��͇,�!�̬L������@.����`@ .�!��4}�� kեҾ���Ư�Zm!��t24u��!�P���DL�NZ!���9�!�m��4��%��-!?!�D�d�r����t���X���/3!����/c���Ug�N��������0�!�DT}H�sq( 99�DdA�J�!�D�"v�J� ߏb�1���3�!�D�/��dPƩƉ]���ꂍ�Q�!�NaF��H��G��hA-P�!�d�����#�U�*��P:&�K�"�!�՜\�
L��E٬L|��5�o!��D�����&Ҿ���>=!�dG�}X�t 5%��9`j��K��!�D�,��0�E͂�T���>;!�d�F~!�3��'�h	s�ڋF�!�dI o��ۑ��*3��!��L�?�!򄏲|�8��S����㞣*�!�$�C���U�E}��#��!�SvSVUY!%F�e��x!�k�p�!�$�.xHXQ䋎�w��Jb��=�!�GQP�P��� ��Y�c�ɻz�!�&,l�� �G�]���H<R�!�D�M�H�)[�� �����;z�!�$�}DDU�fkH?��3��P�!�ܐU�����2h�n� "E�!�ςX̸���=	ͤA�7A5!�$L41�X����lk�=�#O,�!���yTA��QUj$&���B!�ٌ]���2��(9��a���7!�ƕk�� �w�B-�J��!���U���j��m��y��
>�!�$�7��%�!h�8 �:�;�n?�!�&*�<��E�3`���0M]�O�!�\l�  *^�b #��!�dC'K���I3N�D�|t�&cY:,!�ׇH�uKM�<ܘ�'(�A�!�\�~F���ԓT|���!}B!�A	�t�bW�E<D���� t/!�ɕE�h�)"��?��lX�Í�/!�� ��i�J��mx@@��L.��"O��Hd�V�"�U<m�1Y�"O4HR��'���[V�f�h7"OrM8��ʶ5X�J�"��y� �U"O���M�+�\�s��!&�0�zg"O���#��s?L{�Z�%r��AV"O�Dc�aOJ;�@�F"`W�=p"Oةr�N���*Q�a���Z!��[6K�`K@o9�4X�<w�!��.u�
��h��Йh����)!�N��C�������ckĜ!�E�g�v��a��b������'H�!��6
�«S� S.$�����!�$6B��d�3PRΰ�H�#f�!�dA�}hL�i��l��aŚ�.�!�dǷR�(TCbc��ce��8�A�11!�$��@&�9a�C�WL�dCF��v�!򄂭w��mH!��_L�2B��T�!�D�`�8Qq'h��d�R����I�!�!�DK5b������6�}�4�ըXb!��$CxX�nӕy����j�;n�!�dH8�.<zҧZ����;��ǎO�!��Q���q��?C�����E2�!�=Di4��LU�-X֥!Vi�9�!����*i���;?��+%��!�!�DȎ2��pA���(u3�u�d���!�D� ��*س2�!��':�!��P=��H���s%xh�2JI7#e!�90��[�-� �u�'̟'&w!���V�q�-��H�1ih!��0dX���垣9꒔H�! �N!�$�	
�:����Y-b�{�E� A!�Ē�5�|r.W�;$ةل�9*!��ٌ;}��2��ҷ#B R7�$�!�!p.���"WB�u;��!W"O���K�E���N��=1
Pa7"O 4떁�^R�Y2��J&+-h���"O6� p�\�(Q&JE�^-$��B"O���c�-O���c�.P.@����"O�E�a�O�c�]�7�N��p�"O���bg߼'�r� sd��BIȴ"OP��2�F{�)*_��YT"O0��cG�R�"�φ$�~�U"O���É�����J
bB�5"Of�1%�؅0��Mk�GS4B�*U�"O����,��M��C�P�Vxxp"OR��3��p�ٲ�$V�9�J%��"Ob�k��9=�X��w� ^0h3�"O\$���+eF�� �KI@�ZC"O�`#��ߵ |d��0��= ��Dj1"OV���J�o�<�s!�$Q��"O�����[�1V�����^X�"O���T��3&���@]�1XI�&"O�%�",��2F�[�J@�rd�lP�"O�#S
��2mn �2j��C�h�"�"O�paW�#Ui���1�G,-\x��"OL�P��5�p���#�`�7"O|�栒�n��P�o�ZL�"OX9�¯�	̰a'ϊ?s����"OT���P���(#Q�B��l#�"O�<�B#a�9��L ��(����u�<y�Gؑ\�@P���)�$]Hp�m�<!rǺL�0���	�M�|�W�e�<���4u9���K��\i��&D�� �ɚP��`�pAC�6
\v�"OL$����(W�@�H��/H�к"O�x���@z~a*�h؋;���a"O\���[d�ЉS��b���"OX$��&GJѡpL�6r��h8�"O�$
���tϪx�)Z�8�q�6"ORt2W)M����2��0."n�Y7"O����;���4��Uz�"OZ��P�?W�:Y0���14c��t"O�Кv,�&~+p\��$C5j��"O�8w*�6�@sĄ�5r1<��B"O����-V�r,0@	<O��I��"OdYc���mf�lIR(��g�<p�"O�%�5^��^�@�I?^�$;�"O�U3�k��)���]�`�Dig"O�i��d �Ll�[� �IxU"O���6��X�(��f�>�2p�"O<����N��W��dw�8�"�d�<Ywar��ʧ �#K��BHOH�<�P�K-K^y" �Ũa�*���`AO�<�@̛+k�������-A��@f$I�<!� �6�MI�e��sPɡ�(@G�<DKD#$Ȧ�	�擀ba�]����Y�<�QJ �:pXg�K�=2h�"&EY�<�0D !$^蜒w��"+CTY����<I2%� M��I�Ԣ,��I��O}�<ykQ=G礡U��,#�x��^v�<���H%v���>1�� d��o�<��'_4O�^���鏂"mL��5�n�<!��$z	��R ��{a��($��U�<�f��<g�&1�@e�
.�`ҕGLG�<��D.'�VXpB��Z�d	C�<�֫�T"śQEҲp�x:u��}�<y1�Ǳ%�2�bI�/yvܐ��k�B�<M�;.l�q�ܦ�Px�GL�t�<�"#B�ƭ-��y`���;� �ȓk($к!����I����"6���S~,�ia� �t14�N�箸��
�`,��ǂ������ H�M��݆� ��gň�^sd�Z��^�%*~0�ȓ>+^M[�J]�)�|�v���U��hNv��%�s�2Lr�~aD��ȓd۔�Q�'4=�<���I5�v ��{.�af�^'j;���@�ش$K�t��,�@�qlPx�R��`�A�>y~A�ȓK�����h�,z����,Z��ͅȓNӾi��h�,o}\Ik�a�?R|���qބ�#�
�j��8�	ѼG�����aj٩���I�a0q��"U��0��f��uP�	�,��$J��A�ȓ;�sE�?v��z��/����'�T���H�"�����V�9�ԭ�ȓ@5�̑��D-���j���n	���ȓ�Z��	#V�r�t�<# ��ȓp�|�S��'0I�0�r͌��Z0��fe��Kp��>[۠����	��x�ȓTǘ��vK��Llvt�5B>D�0:�g�$��P����B�*5i�b:D��򌖼;6�3����*�(��o8D�����*4 �JdN�"E�)8D�����L2Z� ��5��	'���V�5D���F\�<h�K��>m��a��4D��E!H$k�~,SR�L�ba�"�6D�X���|�L
�nK��d�+�l5D�� �Y�IT����Π@&�x:q"O*���H;o�D�Y��� LY��"OƵ1&��6m4��U��'jR(a�"O���=v���o&g"�	q"O숃Qe�$��z�ȓpL@���"O��k�+MWn�S�EM�3VqZ�"O�0��e�>p�.5�FEơ'(`�؄"O����������J�
NF\�A"O�k�G���hx���)^����"Oz*�W2d�V�����X���"OV�Q�KW�-����� �M�~l2"O�%�����$�
�"O��s���q�t�!��F�|�ir"OD��Ǉ�-�	d��5/����"O��0��.���#NG�h;�"O6e�%ʳu��dQ'�C�'��x�f"O2����0D)4,�$��#��M�q"O*LۡHF�x�1��*ҍ1A��3"O4a�`��$t&����
'O0ԈS�"O �j �3b �x�g��*�:�"O��[4��0\l � 	5@hyr�"O���� р�NER� Z��m9t"O<�{0�3���Bp�P�F�Ɲ"�"OP�P����4�B�oi��$"Oh)ك"�+}j�Y��.\`�L�r"O�ig�F�]����aB�Axn0:�"O�����%��]IpAʵ��:��<D�����-\��ó��HI��p�8D��x�!�
O$�(�6��(�`��0�;D��JWj܁<�\���J�6�.�	t":D��{��C�!YR$ǛA��p�6D�h�"c�9���ළ�)@������2D��C�_�p�!
�"®��/D� C��fZ�u�HJ5��(-D�EI&ZN���-�/4ڀ�v1D���&�C1#��jTBG-9kb=J�o0D�+&Hn`&!�0@D?Bf�*C0D���H%z�)�)ys����*D�����E�B�8$Y��A�#��q��%*D��H!i]��m+!��?Yw�-���2D�l��眾#��h�`���J�+$D�h8�f~��.T.������*�!�$ފVv�ո�a��),�o�M�!��
w�T���ЂX��S�K�9�!�$�	�pj�G��Eg��um�[!�dƓC�n�c҃�QI��KR���C�!��ղ?��1S�뇺[����+ƅ	�!�DVX/��d�6D�XmQ#��;l!��'�]��ҝp�p:�'�,,�!�d��6��k2iF�H����FP!�$�2�!P��zk6]���R2%!�W9Rf"ZpO|��'�E��PyrZ�6D\���u���H���y�N��y�F��Ĉ�se@��1��y�.�<N��(�/� n���p$��y�c��t�A�&Pa@1�����ybl۲g����V�_�E�$�����9�y"��i*V@�PC=�i����*�y�E��k豂�W��Ht���y�-	�'W(Y�q�R�&��5��y"AX:_*��Z"�
ĪJ�i���yR�X
�fҁ�ԋw�9X�eM��y"M]:��Y�em,�I;Q����yB�X�I��M��F�=aݞ�� +'�y
� l�ģ�*h�٪%�Q��	��"O. �'쎆 �P���c
�+�px9""O�l�i�#|=�4�[�,:ve�"O�J�OI�+��81���"�D�2"O`�)���Ȱ7�� K7�0�"Ox��孍�>�Y�n�V2�}G"O�@�Jx��e�Ê[L�z�"O���4��yON���K�<&��ځ]� D{��)ǜb�L��0ԭT�Zd�� N/p�!�䖚$�f��掯R���bd��@�!��ܴ{Ш���I� 5��GLT�!�d_/&&��)��j��� ����n+!���d�������G+8E!�Ą$=�6�#�C�N�R��$a�."!�אBl��[�iP��Ȍr�C^�!��K*32.T㰤�yr��Q)�6=�!򤓱KX���M� &PQ��=(�!�>n���@j��Y�48�	�
�!�ʙ�t81�9!{H��'�Q�!�D��h�Kf�
�AB( [Aa�%I�!��SHh�$Y�0;fT�Y�3!��Y�"��lR�,! �5F؜/!�J�l�j��W�.qr��\>6�!�\� �j<TǛ�t����cٞ,q��$�ZI��E�D2[��umM�y��' cV���MJ�5s�؊6�F6�y��҆X���j���64��� 6�۞�y���(�(sFI[�$ܠ�N���x��>>#hC���^���T�I"C��ٟ��?y��D�2�ݫ�f75����F��p�!��՗Q.�y"�oX�F�sgl�!�*^�l`��eR�EL}!��^�}�!�C�Gn��7��<w���͍�"A!��>�NXSu���X��Yp�#D>N!��Tm�fɟº)�#\�A�!�$]*c6�xQF�!TR@��a��{s!�d?N�:� �o5LDp��B�[�!�DP
w	zi���,)3v����<=�!�$"u��Ҫ�m0������~�!��*&���e�;d��R �#'n!�$O:NM��1AKB5`��9p���AY!�X4b��U�p�Y
k��(�o�=<!��ك_K�����">�����-�s#!�䙊��<�D	�4Q��qX��ۍ1{!�ڷg�t�va��FL�U��Ķl�!�G�Uݎt�Hَk��B!�8X#!�d��h�2�f�����P!�D�\���ꐯۘR�\a)tmH�	�!��C�6*`�R�.�����O�!��0��Y�W�J�m��9�R�14h�Oe"�N����)!�S/g�!s�"O���VQ�2�H e�&S ����"O8�6��X���fCRv����"O�T��.G� ��I٥�Z�V���"OV��G��?)F�PkWmݼk�:`"!"O�-�&&M>���vLG@u8UK"O���fW]�4+��G�&a´yQ"O�U��	5-Z�s�N�&O��P�"Oi�R"� l��i��*�U�\q�""O�!B��R�ˆ= 6��#0��Д"O��5*G�L�~���>m� )�"OX@J��V{�M��v���"�"O"4"u��=R���e�bMB��"O���wj����N�&I�DL ��'����i�? �@0U�0ڜTꢍ�D�$�"O:q��mM�VYm�,� C����"O6�y��V.4qf�̸B�N�( "OJ4�eȆ#r�x������HF=A`"O���Ǧqgj�d��;7e{�"O�]�0@�~�Da�te =b4ӆ"O��C��#>te�µ�P�^����0>�P(�F�بCBeJ5�0���F�<тh�))�N��c��U�z�Ey�<� L*zc.�#���&3�Nᙗ�{�<�3��@u�0L˗n��ɶ�|�<IE��C� 
����ag�Hx�<)Bn��E@��R�Y7l\��P�hu�<��� [���fش�DU;QeLt���0=��
�Oؕ���)0Jɫ"+�o�<Aǣ�&�*0�-k��q���u�<���G:ھ ����(U�bD�F�r�<aK�b���j`@E(Z6`H���j�<���]@"F�Y�9
̔�a�c�<1V��o�B��G�q���q!f�[�<Vʞ�"b�L��N, ��9�T�<��b`�)3�$ּpi4������t=!��˧p�:t(pK�^:��p�J:!�K۴�I4��tY�P0&��.#!�W�r��m1 �Vڀ2�`��i!�$ʸ<"�$c'�]�X@. ��	ļP!�d��W��X#�6xty95gZ�|E!�dЄz�p�*�A��#��cd�?:!�Ĝ	g��`0�^2�`���d_�B�!��$/��5��MP�^ˌE��"-!�+/,X`�`�D�����E,!�D�3�L��$,ڢ8��DƘ��!�3ײ�t/���ꠊ$Դz�!���{���-�Dͪ�:2(O=Q���>O���c��บ�j��m�h1"O�q��m����Q��ꀘo��Ł�"O��
�F�?A�(���)�i�N=y�"O�!�� 	PzF��C���	:"O ��W&ޤD�0E37L[8P���0v"O*����/����K��i����"O␡��߷��MAĊ�&\�n1;�"O���ȍ4!$���/rh�H�"O> �P�V�~�<�x1� �0��"O�i:�@ڝ4��!ph�KǬ�ز"O��5E� %d�yn *_�Pd�"O�h1���2��9��Ԥ9��"O�1�bG<;�"�Pb�Δg:��"O0��b���65:��B=�����"O.�CI�y��E������"O����ȈzF�Ap�L��i�X�	u"O!���:!)�s)X.���"O����G�h�a�b;).�-�"O�٧�)n��aJ%t��"O�EX��Nw��	Ɉ4r��e�"O�x3d@�0���Ň]�L�<q����?�S�Iו9^9��_1xҥУOI) g!�D�WD�D��'B��"�b�D	;Fn!��;#��VC��]�0��E��
�!�$�r�	&�Â<���ɧ�Y��!�ą1o*��6�Ӭ-�Jh3�	�Yg!��G�D�����8Q�(�y�n92Q!���+@*
|��F�J��`���[X�O���dy���eM�h@�.�|S!��M�9��`���Аv�� ��	K!�� X���K�?t�@�� ��I*%"Of ���>/�3�A�\�F�J�"O�M٥.L9P�<"�S�ivI�1"O|�����UH�C��T���a�"ON���aCd:  ����Z��	A��{�A�s2�� O�)SmZ͋��=D����I�!��z���\�	ۡM;D�(H!�xJ*t���-�>IђC8D���t���$�V��$�� I(����!D�,�e��,��u{1�ڹT�&B1j D�p)A׀B��tN��}�D�&�#D��H�+�6V����,����n&��4��V�'�:�M'dݔ`k�h�1;�UB	�'�D�qJ��OY�Ӭ�Whi��'`�hR�H\uL�#��=Vx�	P�']�$���;(�I��ɩL֢�`�'Rt�ԯ��8AAhۅH6`i��'����#+�ŉrf�UN>s�'+t���ڛ+
���J��C�@��2[���'�ў�O��������s�
�u��c����'`�2pkí0����	G�BpR�'�V1��/]+k�.mK0�/:h4k
�'?�y+��^8�n��	Q5-�(�	�'C����^=&pu����UyR�S	�'�(
�o�pBҨ2Ԩb��c�'h�8T,��8����W
�,,6@�
�'��|GkA�9����݈P���
�'�ա�IZE,����d
�'mp���� �JǍ��D�P	�'��� �ѧ>��u�Í~R�ݓ�'�xL�G��'g���0��' ��ݘ7���x��˿	ƨ)1�'	b�9Gd���q��!,�*L��'���dغ^Fl��`F������'E�h�����6S� ¤D�4ҘUy
�'�����%�̵��ֱs�2�p�'�A-Ψ3~��ġ��q��:�'�:�b�	�4�C#H�7~Αk�'���	���4ኄ���T<x�y�'���2�
�F��D�s/�
"4�A���yb�D"���OM.7�lpfKܟ�yR�^49�����.}\H)XդE�y�[�*ɠ�Z$@�%����W�yr��:$Ԕ��aN+J@Ը�w��9�y���y
z]ktK_�j�$$yg6�y�
B�ƭ�!F]�b�APG�
�y"`<e��0FK߸F_:����yR �S��
ƀͧT/�0X����y�l�q��ՌۉQ$��
��(�yB���vTz���H�D�H�E���ybI�S*�p�G��=�`Xs�7�y�o5���4"K�:���1,Y<�ybi^�B�����R0f�a$A��y"k�;�X8�A�;~!(�A����y2�^`+z�!��	"v5��ff� �y����������w��Y֪�&�y���Ԡ{��\���Fb��y���#!>`���.�O����֍���y�n�.B"ҭ1��]
4P��a��y�cΊ�R�r�g
�W׈�3��y2�Co0t["�,GL(#���0��=����$��4�u�H32u�ez�$;m!�D��PdZ�f�\�q�夀!S!�� rƀ"��c �P�CD�|"!�� ����P�}Ȣ1�c$�X)$�"O,�h�D�xU,�h�h����x9�"O �	�C��%S#M��LU�d"O�1��� b=&E��?�Ԡ�2"OX0b@�ϵF
q�!M�s	��	T"O�����W�'$���Y��l�Z�"Ol��AG��KPęy%�?о���"O��KEN٭�-Z���b���"OP�Q�DPx��yw�A�PJ�-��"O�,pգ��F�d|��_�S�l 1�"O��*R(���]���ґ9�z|�u�|��'V�D��j���[;J�2b�^�q'!��^��,���Ku����Ă�M!�d$bY�<z�K��q���(�q!�dU�E�v0��*@3&��i��c�!�B2\�-h�I�<?�a�p� -�!�Ĝ�C���B�%����Y�Q�!�$�f��,�$��9&JT%Z6?R�Oz��nG+~n83!�,8��#A"O$�x���6Er�W� �)�"O����v�"cD��k���D"O�i�K3l�����h�B~��"Or�r0K	)H�X�ǘ 6��"O���	ֺN��$B$H̓]��"O�p{�B	5�N=BW�¶2�4h�u�	N>9*�� ��%C���;5�u�@�!D���"��7�!ˢh��(nRl3>D�
�#��%q<)[�n�=t�>��b�:D��i�펷9��	��1A��X�:D�(�w�L�@���Й
�M�SL>D��
dG������d�9;�� ���<D�(���׷q�t˦h�(OvPuM&�����x�%͍�`(���FF�t}
���"Of	�*���Z<� ��4qČ
p"O(�XG2�����Я8���"O8	j1��A�#A�)Gs����"O�dBJ"��ث��E�n5�V"O2���u�05b�e׽�a�w"O&��5�]�Texx䦞�:!RV"O��󄋪7/�QC��� T�FY�e"O�Ce��
^�x�a䋲u�*(�F"O�hR�-��Cr��tL��`=DQX�"O0h����"�R�hU.A.w:P�#"OuI��a|��{D핒ET�)"OLm�n��ZV>a�C�8n�풗"O���*�Qv򔣀-I�K�� "O�����ܯq���ؒ��-.�X)qV"O���  ��SK2�U�y�r�"O`Iq��6w.x� �U	D�2�:b"O���j��V���ӂ�S�t��"OL�� ҙD]$m�g� �hD�p"Od����eJY��FH�z{��1O���T���s���c�B��]C��O8�=E�t7O,U���U�<�"eK��	]*ЛD"OL��3+92M��[D��5pP�l�$"O@�xr�TR�w�,'X�AE"O�Dy�!ڛX���qi�]�&��&"O2�hG��+*Y��
L*F�<�B"O|�f�хx�6��%��.vVP��"O��À@��f�tU�ehI7p������F>�5�<`����W�M?8�&IW9D�B�%	����£���EId(�e�2D�Wd �/Sت�D�:a���0D���V��0*U��nM�"V��*<D�� &�k�O~ch��Ԥ	���L�"O,ٻC��G���0�+�&�3�"O�i��[G�ZA��"�7��P���'U�O�}�EKDpc�%�Q��C��!>l*,��L���0���*6�y+&$�2+L��ȓY,�P�* 抬�􄇗&�����8Ҥ��d��Ij&t��?s��Q��EL��6�1(��t�5��c�l �ȓ;/� ���\@�=p��+8ߚ���Q� i��-I�Qƚ����(#�x؇ȓ6b�x��J�@I���g������<(�祚�
^.TaR`�6D����UST��F�O�&[��6���0ݘ���u�ބ+���-Am�
V(K� �[�����̀�h�;�L+�d�ȓ6�z�aA��-O!�Q�ȓ+����t��b`�X� ���i��	� �B�5sf�&�ŎU�fh�ȓx ����;۠��*��[��U��9���cx<4%��K�\0��(؀�H�ǔ$*d5
�郝V�̉�ȓW�F�z��[ pEd��/QkH�t��(�d�gdV?0���p/_-=Ld��Sz��Q�N�,������$��?y���~��bj�,t
�挲[ �Ѱ�/�K�<�1'Ю4��<�,R+!~����~�<�৉57��D�w�K(8������W~�<A��;!؈I�v)��LS2�ð@`�<���� $�Q�E�o��u+�`�^�<!w�O�r�68hu��(�R|�sD\U�<��o�'r���!�jˡ8��e�&��H�{y��O���Y5[R�B��Uw<��'����Ś?�.�� ���&�,*�'l2�9s�<z�A0�	���j�'.p`bn�B��ь	�� m��'������ǥ"n���M��	�'��A!D�@.& 0͞=n�6�	�'�dh�A��T(dKϬ;�(�L>q���?q�'DZ�����V��ة���x{ָ�ȓb�0@�í��9�� `6Ĕ�> ���z̫��L�Ov�=��o?1Z��E{��O�����ŵ���;�h�v#��#�'���a�GU��`�Ri�w
���	�'�T;�D˄&ܢl�R��&z����	�'a���G��6W@H	CF��P���'��d��:4N$�����w��Y��'7��0���-(le��_�qZ�'� X3�֦a�����d��^�"���r�)�T�����Y�Z>��� ����y��Ʒtl���G^��9��Y�y�C��t�r=
g�T8j`������y���J;�ٻ���6�Xl� ���yB��;b���J�R42_�]0���:�y��2��<)�a>3�F�KW�	��y2$J&A�@pC��3�hu"� ��yR��#L����^'d�հ�װ�y2f�4*,P	)�a=$���y��^�y"dɱdd���'P@�6#�yҤ��Q*���冎�}�(QHW��yb�"_e� ���,ec
��3�yR䀫|Q��P2�ݎP�vx��V>�yȍ4�����JZ`����N�y"kQ#P�b�ç�J�C�z�8�c�<�y�×�	:�<r���r�Z!郬���y
� f�WB=����&nٔLT���"O�9 ��[�n�8T*���:]�ZE"OLP"�V�Q����M�,ޕ�"O��cL]��&$��A�'(,�8�2"O>�"��I�-jqx�g�9�jQ"O����H	�P�� �@��'r3D�4"O��燘L�E1`L˒Uv���"O����+I�>���r��]h%��"O0�Yg$Y&,@t��ԩ��6`*��"OБ�hT43*���gC�d���f"O<�F3wkН3���c�xă�"OR�aD�ԋ2CdT�U��LtH4"O"�*"#�9�ꀯڅ0b�E["O��X��i�዇.�#([<���"O� ХI�J4��1�1Jh��W"O1�S%�(cUn��I.�L�Q"O4X��T�h9)�\�O��"O��S�ċ3���$�#m�݈�"O|���O��՘�Ň K�`�h�"Oz-��_�q�"��������"ObԹ������׬ؽ+q�h��"O`�x�d�n�^�{�ID�r���s�"O���d�����a��7U-0 x"Ou�a 
�@���G�	#*��"O�0fb��>~�)jf̏pT��D"O���:��3EX5##޽aW�'n��{�j�P�6�1���.�B�|��!�L=��`�FI�K$�B�IT�[��� 3�(�'�G�]i`B�I�82=:�Ƶ6��!AN ��'��'$���q<\������:3��3?�B�	���\9��҆{��p	E�V�!��B�	cz>XZ!D�>gCn4�A,W�-n�C䉝LaC���mĈ=�07o�C�	!� )���̹<�& 2�h�QʢC�*/�fYȁ埅a��-[&�
�HB�I�3*,u�m�
Me�����Ǉw�B�=1ç	�����_�o��P�)ݕ*J��ȓ*�.@��$\�Q��;��]�@yꄅȓd�����׮.����S�Nؼ��l�'�I� ��2E�
u�+�J�
���'��૧-� ��ģT�[�<�%��':b�1B�� 7N�	���R9�0�
�';�]Q��N�����+g
���'��=���h���1M<f>������-�Of2%d�[��Eb0�&?�L��1"O(�it�y4�-��(N)lA$8"�'��ւVC �\�C���vر�L0D�LC�� )};6ahf��<�2�g1D���"��^��;S�JO�H��V&$D���c�X?K�#F��@��2�#D��hTE����;��B~ }z�D#D��[��_�1�����^8����"D�Ljt�
b���rK�|[8�)B�;��8�O ���jJ�k���S��W� ���Q�'��'�az"3��ESԯ�1S�R�@w���y�o<>fʡS����)�V@J��y2�Z`B�Z�mZ��rh��"���y�ė&n>�E��$bZ��%녅��x"�>|.�eçA�}FpY0d� ?�!���&�	S�.).�@+Xn��2?O�Yɑ E�/*��8`�է<{�Ԃ�"O�4ò[u�d�G�.jd��(v"O�\�tM��h�NI � �+��XJV"O� ^���Y�L'
ͦ[\(@9q�'Wў"~
�&��c��qJAf�]��`����>��O��L��}�RA�D�B���R��'�1O��qSaN�U6�)���l�>�""OҌ��߲�`YjM�Y�@ A�"OT����"R��y�C�:q
H¢"O��g�<@���l� \ ���"O~��U	Ҫ ����ȲD�<Br"O�1����h��!S��V�@�;�O<�hb�:�X�Jc�B!#�a���)D�؋EbL�_���#�J� D�81X���Ov�=E�4� ��@ȓ"��g���1�#[�ўD���),�� �@�,V4 a iB�I7P0�(�%�� )BXYb�Nrc�C�ɤ\Ƕ���bK�Y?$��0��\|B�	48Ȓ$&�"��ӆ��H�^�O��=�}z��5D~1����zL,R#!�c����<�S�Q&H�b�J��<�Py�v�@Z�<��.�U����Ƿ[�t|��PA�<����^xd��Ǯ Ը�Lz�<I@��s���۰	ݾ[�N��s��o�<і��;�v4��$E]܈�� �i�<��猐U�FU��j�$g?��GQb�y����y� |���D!�7
W�3"A��yB��B4�]�4C�	U���!����y�IO5egXT��)�q�Jx�(���y��
XL��
f�Z$�	�㗗�y҄W3:��;���?��Z�JX1�y��]Vx�+v�!C�2�#�$�.�y2LA���S$��J(��"C
�����?�S�O�B���dӈ���I�'0!r\�K>1�����W�8p��!A5*���+3nD�{�	S�'V�	j~�AD��'��6^��9j�(4��7�O����ʵ@��P��]82��ٶ"ON��rÆ>.��)b�#)��Uу"O,]!��ҧ.�3���:���"O<�;���"4.|�I0B�lNrT�q"O����/���s
��) T���$'LO%`��Ȟ9gnY0�m:(!�q�'Z�	E��!@���02�����Õ*�jB�	~�nT���Q�:"<h�de�3Z��C����)f�U��$�xd��C�I���И���//��*���1+L�O�=�}��e��v=���4N��FH�;EQL�<�F)�̓F�Y��
��a��^�	cy"��<Auh�>kk,!��R:x
z�zĪ�u�<���I(b��z���=�vY I h�<��IL�D�rТ�C� *^�8c��b�<	����F��seh�;n=�U �e�<�1���{��#:%6H��Q�Q^�<���O*;^e4��7f���P�/LW�<�Pn���]��*dJ��fT�'z?���J�3P�4�b���q53A�5D��֭�9@zU�������H0D�Ԛ�Gȗ]X��1H"�V����-D��EB�$9| `r�	dv��+Wf)D�ҰMΙ<���%N�.=ߦ5��&D�����f%*��ϡ
��	y�.)D�KĄ̱)�q�G�Z���%R�'$��s���S1X-RB"W�c�B@8G��:"VxC�I3���r�! 
]z�d�ۆ9�>�=Ókgt(�d['�6�*7	�W?��ȓC2���[X�H`�0��,~g@��[�JA�B�V��%�E�)pw*���S�? ��eN5a��FYp�k"O�╉�3~P�D���<`bMqC"O�`�5bNt:�Ț�j�6R�-�3"O��8���2�$	B�V�.=<Aa�"O��s�����h�	ڪy��"O�ca��?`�$1Q7F+'/b���"OZ�����6>� 1ж���l8k�"O�)��c�V�x�#^�G� ���"O2���
�[P�A�ǌ�c�"O�ܰ�Nޑb�uX� �(��B�"O��AG�L�N�<�h�/�'h��� "OV�y�^�0^h���(ձ4�Ŋ�"O@��s ��&��+���H8�P"On�U	����P��V#�A� "O
���	��J�T9"f���0|�`4"O8ͻ�g^5-���!������X�"ON��� �) ���j�	Z�r%с"ON�@�FJ8.��J�U
q���"O ��p �;HK��t�B `��9�D"O&���=�V�S�G<>��ͺ�"O��Z�)ɋ4%\Idj���Rб"O�a���&i�� �o�z�,PQ�"O���G��gX�L@���J�l �W"O�Eˡ��8D��Q�����ʁ"O`��vO�<HH�m2���w"Olpk����+"��b-J�i54�"O����@��2�j�ړ!�sD"O�1X�Ѫ�A8b��x��""Or�UGؘ_jj��g��⁣R�y���,���7Ǹ;�MAՆ 7�y�i�="�:ӧ5����O���yB"��By�r@T�=M �j7�y���Q�( FgX�-c��:a�֑�y��6PW���)��0�0i�3�y�$D=�a�V��5KXd"ѡ�<�yr�V��\"�]X�(�˵!��y��W��*G�ͦz�VQ�$�șE<!��E-�rŌ��0e;g)Y8B!�$��jM2�G\�K���:q��"3!�$�(��Pc��G->���8ҥS;+-!���1}h}��Ö5�xM�B�U�!�d�z��CR$ښb�*�11�Ք�!��Ş��0���tc��@H� 4!�O;0J�� C�n�8ʇ��C!�䏂e�����m5&%k�&32!��S{JHB��D�M�����V�!�[�F���&թx�P�C�1!�$T�$'^��A�ň\� �s!��?$!�D��u5<�JG���qCp��cʤ8!��%hK&I.d�TI@�E g7!�dɰ@*��[�(����_�X(!�DΩ����@���J
(��gN�c�!��3딙�ѣY�2�"bf��6%4!�J�4�9H&�ۚ����F�J#U!��Rx����HM��h�!��5V!�Y�^;��;��g���k����!�K� dA��ėY�
�1��R|�!�ė�`�<u�נ�y��ђ��~�!��_���%��0�	J"�U�!���6��-�b�{��85A
�j�!�dU�G2��z�l��ǌ1	R �;w!�DE&~/��
3a��J�`�,εS!�$T3rƸc�Вx������#W�!�C�64h�L
 b\h`/Ư}�!�� `�ۡ�L16������Sl��6"O>HA�A24�)Xt�ڄ\�(�0"O�x��Z YT��6LL8�6X��"O�uS"P�F����]�bS\)�a"Od8k1�@�{f<YG#�\e�Y�e"Or��v�
3E�$d�P�,1dtX�"OD��LLצ��@F�C,�t�4"Oʈc	�� �-v�и6�lPcc"O0U[���j&y��c��J����"O�<�p�ݞJ/��bCaɑo��0�"O� #%�S�L�5��6>�X7"O�hq`+��,����D�^�j�"Od�3�((�:���3-��9D"O�I2a�6C�. ڤM��oN�{Q"O$5����:��Rvnb��8i�"Oƈ@v�ö.�� �)�MP�?D��0$#<3�.�y�JV�L���>D���p	�7pG�xq�Oe�DB��<D���#�Ѱh����w�[�VR�l��/D��5H�Bo -H���x��O+D��Э�=l���T��#`N���+D�jQ��)LQԨ	��]�D#'D�Ts�! �j�*���]��h��(D���'�'_{:�-��Ԭ*D�'D��0�	��	�ݘ���P$�t�E�#D���D��(�f�K��>#��t�=D��r��c#t�82h7ԀdCa!<D��
bM�8hdZr�ܚk�j083�-D� g
 �nC$�:d�Z�i�<ԓb�,D���5K�!	��4�ř� �rȶ�+D��ГŒ��L1+ ��.�n\1b�)D����x	{��"c��HcH%D�pbwǗ�w�2t��'���R�>D�����T���`�%�_s���D;D��*���-v���J� ?H �h��3D�hز�"d�
��r�
v�葂p�2D�$��-F(�*a
@��cN��5(;D��`��5}@8��
H6c~,�4�>D���h��V�^l+���s����H<D���
5"D�[�M�_ޙkvg$D�x�HC�P�=�DB�$=޲�j"D�#��<\ĳ��N*	5d�z�B?D��ꤩ�4"��u�MQo<=@�8D�d� M��8q��f8q1�G7D���e�6�(ف�J4w���"��6D����! �A��a2S���v�J� !D�|��(JX�H�À��\C2��!�>D�LH�:	5DQKr�O�7�D�#v�'D��k��ݕTN�aa
�	�(�9F@1D��`F϶� �� �f�Q�B-D�H�v-�_�<$�1�@�(�p͡D)D��S�P�/��y9�o��3��41);D��+�@�Z�ec���A�d�)��<D�����V��O\��2t�g&D���t�2��U:q,�$C�>劗`2D�H��XlC"͸�˝�-�9�a-D�����2�����_��У�J'D�\�a�*E��:2�*n� 5Hd#D�$�d
2 ����̡�J	�q� D�x���#u��c����$���"@�1D�� ���}/�	��ήIނ��$-%D�$1B�I0�� cK�AцЫ��(D���Ƨ=w�p�%�E�m����N'D���3�4'8��'�L��1�$D�� �H�j�K�Q��^�5�D��"O!��jِ�����
d���"O��as�L.&�T��b�0��"Op��B_	��e��C� |����"OJ�[T
��`����y�����"O��:�N��o}��z�"_�`�� "Ot�{r)�O���a��]�����"OPͣ�l��I��م�6�b�p"O��y��K$�߆m�Zi��"O�������0���@���0�"O5��t��!S�&������'�4`��&ԧI��
�`T+Nx�9��'�ک�V@M�'����H�x�z�'j�!���	������ݓV' ���'Ҭ�j����\�=zt酎K�R	;�'�\����	��ezc�	�>�4��'�(ԮF,I�L9#jV�:;R�j�'| �vk��4bB���3c��X�'-`0{ECu��@bh	.Wξ`:�':yZ���58��@�Y&��	�'���kC%L�[N>�k��R�{�n���'���kL�-��u�3h�1D��+	�'H"eR�Ѕ>�D��Rń�6��)��'�ލqe^�+F��H��T����'#���c�O�u��,�Pʔ=��U�
�'�>�B�n�f��IQ� <q�
�'�а @��
���
�Q����'�F�kŅR�5�~�y�	���b��'��(�Wg�?\�$�"ra�Ҡ���'�D����>'����k�a`0�'>2\���[�4a��A$DJ>{L[�'�}�pG�W0�����ե_sx%�'\�z�g�Z/L�04��"T3��r�'��
s�\�"!�	���8Qb��!	�'IVZD�tߊx( BΎO�>x��'RxA@���]���G�I�]��'jP������ĕ[�/IF�r�'�Гƅ-zJ`h��N+=�~P��'րP�F풋,����D�;_+X��'|�=Kg#�<�xTr)T�Ic�:�'����tM'lJ|� J�H�����'2x�*�V+�T��h>4r���'�&t�L
�	$R��5���;!�'v@)��(t|����N�8)h8�'���3`9��l.	�CXf�@�'/B�c��$I^���N�><�b�'�ʥ`� �0�vh�s)Z�0:t�A�'�L��%S�0H��2f)�.2�h��'����"Ɂ2uB����h�8.a�T��'��1���B*jӬH��"��"�d�(
�'�x����ҏ8Q�P['�»,��	r�'ː�R� ֙nJ	����$�#�'#`���0|�L���] UZ���'��,iu�F�S���')6���YD�<�b"���7*�A�^��bjWu�<Y�C�t����v��{����V�II�<q3Ʉ�-��șRK�u(Ő�,�C�<y�b�.V�i����H*�)
gJ}�<Y��N>eLԥ�s�Y�}�4�����@�<!��2@n�J��� kB����LR�<� B٠2!�y萏5��m�%*T���Q	]�k�,�5���`�h�aA9�1�O d�a@	pX�Mk�@�]�ҕ���'C �n
;�Vܙw唴 �|y��?(fB�)� �Q���ѵ�>�����p���4�'ﮭ����P�����A���;��8|(}��Y��4)Dn�sѶ�ˤ/�,lb�M�ȓ �q��G�ݱ��R�.����ȓC��a7iI,�vD����B�I<�H��	�Th�@��[�zֺ�����B�<�#ǟh�R�9���k3�B䉿>�EbU!�S�8���@1;����$�"���f=�e�K�%M���16`��p��bH���*�'����fnN2+���=�����$�P?h�@��/�R�j����yB+O�
&���&(��qA�斛�y�G���{�!�*K��IP��V0�y�g�H~�!�JQ�e�a`�$�y"N��2�Pz#�_�R`��.���'�ў��,uآ
�w�d�S�]*3�
�"O��hRQ���2��Y4~zXr��?}�)��3�����O;%p9Q�@��C� v�$2`F���X�kv�߿y��І�I_��R��L�A�P�Ag.������d'�D��xUI�M���2�Ĕ4fQ<�5�9D�x�$�����r5��B�ޕXB�I�vь�.�����	��[�j�pB�	'<�R�3���7{�5��K�~V�܇�I�HIt���iUer����G�-r�>B䉱e�A�!c��B`�[�܇$<B� kn�ءo�<AT)�'G�Zo@B��If��E�r��-ѬP8"<ϓ�:e���+��T0���e�VՇ�@k�iZcb�4Y���U�E?:�rm�ְ?�2IF�zHZ%����t�N�c���<�N|j!ҟ4Xq�g/E eJ�)�c�N�<�2h��/��������,�S+c�<aU���	��y�+^�h�x��\�<!���[FL���ɧ?���8&�U���7�Ӻk!
�Z
:�H7�9�\B�d�R�<����U��m��L�?\�ʂ��P�<�4B�.>j<� m�9|�y�P�<Y�K��2�m�tƜQtf�Mh<Y�� 7L\�y5&Z�ˌ��eG �y�(�>BR�p2L��̤²����<A�d��[MlI�V�"0E�){E!�$9߾-�S��)f�*p�Dlc�'pf�Dy�dƹ��	'o2��Q�`�� �,��ùc?�B�	,+&y��
¿;��bf�\"<qa�	]y2�D6X6z�ш�	C!ۤ	V6�y2̖�l2V�R(�$��t���y��]`�p�ku��<֢Da�Q��y�*F!vj=#�gL,>xUbG��7�Ov�=�O\�@�W�G�)����kK�fi���'/��aT�D�4��8c�_[� 
�'��H%���Bbʀ�BuT�c�O�=E�b	�h�6�悈 nv�3eJ:�~b�'3�dy�*P��Ճ�m�0�\)�J<q�
��I�	�x���۸�Z s"$�zE��$*���e�W�1��r/��4��`�f %�a��#~�%� �Jrl�d'˲bs���OP�<Y&�#LV��+Uɺ`A��\I�'�ў�oq���("��� p�Y-'��ԇ�^иS�`ߩ����ħ̡��l����a5�ݫ%�F	�7gY��0�ȓ7ly�2g֒T��E�0AZD�b���_�MR|B���6zl�#�M�d ���Fd���@�ұ 8,��H�-��>Q����� ���DmO�@�T0�MGt�PY�"Oj�14#>�ARP�e�4���>	)O�R��Y��Jvl�m�D���
H#H�(Q�C�?D�Ij^*"1�T0ISP��DC�}��C�	.4B�y�̎�{���۔@�>k��C䉔[Ŏ��� J��fAK�'(����>��ʏ�a�Jaq�LM�/��l�t�V@���'��	�<1��Q���cXZ7|���D~�<���6hʴ9uO���U��(�v��?�J|��&�6yl9���!"�-j2��z�<����%�8�R����j��P��i�R�<�B(F:�X�ŤƑ�M�O�<�!@��<�Y�b�)jJ(�Ј�N~��'� �y�O;,ڔa�cd~�@	���d�o�Zd*���M����ǳ(�!�$�~���#�ʰ����ߙo?!��:v�L�Z� ��$tę
c�U[��.�Ot0BbN!�N#!��?���I��iў"~nZ�thE��b9p-��i�+0"?)��鞓F���)�+�
iu� �ԡ�D3�O��B(�`�2�1�&�F����"O�!�(�
B�H�f�3rJ� �!�D]�B��X�1	D4�>���!
�2�1O��	�����'���HP�&J:T�f�0@��%�0?9-Oy��H��"6�e���-Q9��9$�iUd����dퟱO��$�B�������=��-��D!�䋄/>2)i�
X2z���J�l]!򄎱-P����A�#}�A�P��!\a}r�AyB)�F���6)��}������hO����$�]�P�
q�����W��4e�D1�S�S8>�&0tނ\hp��2`\)�*c���I?TN��2 3�eQ��<�7�͉��I���x�%�$�p��'Sr��Vn���p=��}"�S;I�Q; GŒR&�i�f��-�y�P�Z���M��E�R�:wA8�y���	��HD�T�r�D�F�N-�yB�]̠��գ�p�2���-��y�JϠ?Z�P3PO��a�X�1����y2Á%	�!�5��<E1D1��/͊�y��X�2��MCv�&��衎W�y�Ì�fA~�cEX�PJ|�!��y�!'
M�0̔�{��4x1j.�yB��8W<&���'��<[����^�y�����T*e	�~9��P����yRM�yd5��(�7z�!hw����y��O�_��X��[�����v�Ѓ�yB�#�J����̥�T@���y��<t���يj,�c �7�y�\%���B��,ꑏO��y��Y���Y�`����Va��ʡ�yb	Jf�8�f�h�ʴ`�]�y�'͟-�H�����*������y�'�5K�=���X��F$	�y҈P�lS�x�$HT�]i,@�5j�y�',0^�%�i��S��e��8�y���w���� yz~��1����yR��'I]�TkփX�k�5[��=�y��	O�(�p`�;]���#��C��y�
{���3��O�T��2�
�y��o�����҇^9�ȱ��y��F=<]	0��3P��5[�1�y�
�-�ʁ���H�}t�B�	�y��6{7��U&���p�lT��y� ��e|���`�=��$�����y
� (��dE�9�>Qc�2g��� �"Oʄ�s�O9�ʐQ�!Q�u�zu�r"O�(xlۺ&I\�U�0ٔ��"O8��c��VҰAkр��&�4��"O��#�B�L�i�O,}�4��"O������yhZr�MI�V�&"O���1���a$�r1���t"Ol��C�<����fe�=���@�"O&8�T�T�7Е��M q�h ��"O��RB<J����S�B�v�00�"O�в蕟o��$���Rüi:W"O$���O-?i�1 
�&�,X�F"OJՋG�I�r�|� M�IL���"O���U���j�­Q�M	�iB�5C�'����a�,�����T9,,j�)�C:���'��Ps��{��D�!$4��X
�'�PK�n�{�R0H���	�@��
�'��cF!�W�6$y�eܞ	x���'X��`0h�,H�H -�rnf�`�'�&,SV��?e�"�*�ޙsa��'9��xAŇ�2� ���qU�Q��'��1�3
47��SH�(:q� P�'0������]��(�")�?�p50�'�ݻ�o[�Lc����ʢ(?���'�n���+%!����m��vfj�a�'�֤�E�?
ʠ�I
QvU�l�'���!�b]��B����/n�F�a�'�������m��]ڲʉe�d��'4�eۆ�Z,yF��reħw��s�'�R�k�	ىAð�@"�ڲ�`���'攉�@�j���G�� z�'(ɩe̟�Q#�Ջ�'�y�z�s	�'�ăS��&v����+�èx*�'�֡�B#lӦ�1���"�J�'�0�zQi\�^�@is�v�6���'P�PIP$�Q���Ctϖ:���H�'!�E�r%W��n��#�x��4��'�Ӗ`�
O�d�kR��)D�dUH�'\T9�0�G�t�z(0Q��'6`�q�'��14A�1�|��,��8<*�'��mk`�S�p>=��l >�P��'#rI�'GK�V��C3ꀗYz�	�'x��P�Hq\�9rĞ�Xz��
�'&Vy��8re\�F�L ]��R	�'��M U�4,���`�GB�J\���'�2�3lޭd4�"����Ɠ�y́�j�yfu�t���yR!0{1Ԝ�F�[�D�DÞs
�'��<��h��a\"|�� [�yr
�'��C��_�ʰ�A��}c�L�	�'nFE�3C��C4Bm6�W�u�^�H�'˸j���8Z�h�F):����'oXR6�J�_�
�ɤ�N&8{�'X�d[�Տ6X��JF;F����'l�!�+N�Z�܉0�[`,�C�'8�􏎀�0(��W
�b9��'�~!���	����d�V�!���	�'?�h�"�7=�a�S�֭T5�I��'D�ШR�z<�A�''Y�C��x;�'�5���%�)�
��J�X̐�':̔���Б#��P���t��ѫ�'�������0��!�P�Zd�u��'�D!V�*w����7D����'�l��Dʖ])ԅa��Ҡ	�&��	��� z�ǉe	*] !X�p��S�"O�q�d�5޸Epb�9-��a�"O!��KD�FT^e� ��W��\@3"O0X�6L�'H�x����.�x�"O��ju��=c���{�q�J�P�"O��
!	�r��@5	˫ΆɀU"Oʝ1f��9���jL?I����"O��Q�	�>���w.΍��4�"O�u�`����.�a��� �<�`a"O�L8���%l:m3 (��
d(�ї"O.=����,S8�(�j^�mXD�0"Od���r�I{��1; �Q"O&��E�Y�,��=�ǧ�)i}4�{�"O~��k�<󰸣R�FZ<�R�"O�|�ϸ6��������9�1"O6�� �^�U��(��H�V��""O8��Qe�����"B�J��%�"O~,�E`ξ�@hv�Ġ�|�I7"O��qF��
a���2���C�`\;U"O6���NШx`�����Zd���"Oj(��O�U�f8L�.I!�P�<ɇ��6����%m-y��1g�z�<��ɔ,b�̻�ņT�t#�v����9��{�� �7*����EC�d�!!��y��4X�%r��
�*���Xf�֨-i�'���p6֩��Ϙ'�|��Ĕ99��bKN�Ai	�,/<�c&�Ŭ����Eڣ����3?�ܸ8�(�[\�52	��l��y�!��g�x�	�BtGx��l�8 ɳC>X�"�pe2�
.4~tt����L���N�I~!��1w�*%�
�`q��]�Jg�C�I���ʽ0ь�U}֍�d�i�q���9�4k��(�0 �.��dB���g�V�<q$�����[=7oP�Iu�J�6��t�`bQ� &��C��U�R��(A���"�%�,Q�;S\��G���� �'��a��3�1����ZUR9�a(�p�*�N�/j�M9g��_�8�'`�(���J�t`s� }��蓶M��eǘ�ҦkJ�n8Q�H0�ɂ#-9��-Z/o���MV�<߉O�!Bg�9[��D:�R�,RT�'!��"�fS4�bm��I&n�BN�B�`p���4 Tp��"��LJ��%jo��I�)�5r�0 1iۣQXz����R"Q�p�� E6^�P �' ��;d��= �nѱ���?Z�)�i����$V/>nl���
> )�_}H�y��P�K���YD&��
06���N����D��iV��Po��M�����W�!�AٵnUB�İU#��S�t�:Ђ�^�R�'���F��{�!���OLH&�02_�FxR��=A��s�j�7,�����D	gf,�aįrt�qA���~B�ޑ)j�3��K��XHU�r�d�DY(?�>�Y`�ͥ0�RY1�떟HC����c��O��(��8B��dFЪ2���c���<=zuE� u��=�ȓ��H�
L�S�Τ[�凾B͜Ml��V��7�٘v����GHٲ��%��(�X?y�Eǿ@Ϟ�0z眭 %f8O-�%���/L����`�h�C�k�����k��W4/��M� @�
���H�G�.zp]��|� �O����+E�߸��	Cg� ��L~@��U��Zt��2��.��Æ@�	vd�}B�Ɠ�l�
Y[�C\0P\nhA%C� h0���&:���Ē�,k(�蔣�Z���Cf��k�&��2�C�J14q��J	�0d�1�_>���ŗ�"�Ԍ��X�lg��l��M�Wgɽ=ۈ �f�<D��)��Q�q�2��F �-�d�A�S�}"�BhV��i",�!M����ҍC2L���5�:M���_(�"��Q I "����ߨ�.���`��'��Mcj��j�#�Juy���ƚoJ�]k�8���7؀���Bm�3}"�
�0���SG��r0,p@��r3$d;�%��h��PSS�:v�  O~SD�C���ȓMؐdłD9�M��IAHPjĎ��?݀��d��B�5�G I���ɳLQTq���$ې^}�(�$*�=�eieW>�S���%}�<[�U��5il�6�q��(�,�Մ34�h2��W�H�����LB%�t�X��vI�4�N��8d2AAȧ1��#I>9a��&3��ϧ#��m�U$��. �"PAT�D���/�b�g@�R�^$c2JiC8u�-T�	�mI�A��<�V�3�	,ND����IF�	s���"sK�@���B�j�*\iL��P�	�G��q��W"d,�z$	�?Y8t��żCF;q�X�J��b���8V��OH<��� �:b�ꀈ*DϿMʼ�D�%y.4�.�*!G��ˤ��N�2����i9?)��� ź�y����lqp5��d8��F&A����Ŝ�P��HD�r�֥��B�&y�-���K�N|�3f��g��Q�@~8��rB%M�(�Vq"I�tz�`#�.}b�����(C�ƞ]~��� &��A���>>��Di�Ծ��XC�Å0��=�`,�=�L�;�RY�ƌA3
�Q���M L�ÍE��I>�6(���+ޒ!H���O��C ���yG�SX�=�b�� �<�֍İ�Px�	ͭ���qF�X]�8$LC�Mς�Z��=e4 ��E��B��lH�����CA�Y����͐n���n������7Ob�y��K�i�Of}�vgJ5EL� �o�tU�wlV7kq�|��ŏ	���n7<Ol�B��&6`�ax��L�Q4�>Ѱ� 82�0�( �DAvh q0� ZF�P(��L9�����}{n=�b�_C�<�S΂5��,�"�,Xt���dF�= �(�O�l�q�gwD�I�����B�S����B�@��LӰAπ
�E*��� d�!�P����`w�X�e&�kf.ψ �Ј���q��ݤO9��c���J'>�y��P���pw2����<ۺ$��qu6�	Óx�&U�Gr�b�oSYhj�x�ʓ6YiV���d�(�:U��n�]9r��[�,����ɖ pن�	:
�&9P�� ]�$�iW��	vq�p*�MA�"9m��$��d\l��ē@P�XT*$Z�}C���")�>i��GJO
I) �(Zu�`���D�8<S�Y�#^�l|Ȭ�b��y�ɔ�n� �+A.��f�" vE��FÆ��?��ER6���Mc��>�6�DS�L3.ڹ�3��ib�C�#zۖe�SaP�2��T��ə�@9���٧>9c�L~���9d�9Ol$�4%�
����k�$D�1A��'����I��fF���Q`ӗ+/>Lc�ɹ�z-�2��!dpH�BCt<�u�8n�RC2Ԯ'B,�U�FkyRLIQ�>� ��V
�nm�T�*SȄ�(��)�,���dJ�)�B�8ą�,V%!��߾%�`,{$H��Y��KD"F���#��ǱB�ġ��{�N0J$�����)�z�d���S�E�?�b�3sN�nO������/����7OD5y�P����&��`�ӧ5�J(`��	�6]����%c ez3�'�,�A���^(b�#c�H^�ys���R'T��%bW:1��AE�5t�"�yD���E#1��!);6�Z0,��hF~��	�'c��(��a	S���=D�p���'#^iXSș�{�=��+O72�^�HD��2���>�ʵʐ�o.8�G#0�ԽY��$D��
`�+4y6��ԩ\'lhb�$E-b�j�'9M��U�v��"wC\�O�0��D�xBb�?9X`�a��
i���F+ބ�p?�g���/� �qb^�~�d�D�WO'Z�0�AX1+����gɖJ�x���0Ӫ��Ҍ]��VfِQ.Q�t!S��)��=+��NP�M���jU�8Eh����Ok B�ɶ+"��#$��h��8��4��I!P��Y�� �����h��R4�W�vL��s�R�VB�L�r"ONe�ȏ�G���B��U3���re�4}�ƅ*d��٥�(��DQ��nt����K��=�/řuh��Ѽ	�`�i��Y>(�|�q�; ̈�BC�'+!�D��^���TDA���M���%�!�_4te���Ό*�J�r%��>T�!�dӚd�"���Ɏ�g/
�I�H�!�Ĝ�/2���)��Qm�i��7Qv!�D�M��uД�ϩ;Q���VbA�ac!��Ȟ|�6��.3+j�Q⊷Y!�$>� ��sg�>s��� ��!Z!�dF&�:I�����[����ѲHH!�B�O����w�_�]��HX-O�!�!�G4$Z��&g��Vt랠#!�D.@<P��a 0hxl�fK�(f!�$��,��2�PMZ,����['S!�D�-�� JRh�sD��h�^�(N!��!	*���	��-�dj�5:!�$A=w�TA�cq,a�N�V!��S�.�pQ���=fP�S�&H�!�d]�L[~��)�0g4,s��޲&�!�D	�g�6�6.ځ7�9hע��"�!�$݇=�88� �
2z� �bʄLc!�� d��GV�����ɸ|~��"O��bÇ����.ګK4��"OڕЅ�H-
���l��}�""OB�� M���{b��
Q��TX�"O�݉S?Ԩ����E�WM2�"O���%~p��X�/X�T���c"Oz�*](�����e;AKǮ[7!��G�A���D<�yU�(Y:!�D�[�$Z�+ь��F��g�!�D"\�{f,�+3��=>�!�D.������٘�|5W�3[�!�D\7$�M�@KV%3�X�$��k]!�$)J�� 
�K�}���{��ٙvo!�d������K��9(�#q�̀SJ!�D�-Y>���<DQB�ǐ�+8!�T�:�b gE�g�!s'皪G!�$�(.��Hҥ؛���af�;/!�
91Kv����3=2b�`��<=r!�d��g����|!|y؂�X�!�D�2&��1��0L���*$e�!���wl岔�^����:�!򄞊%��S�I�<�����!�ęK�*�z�'[��|�ŉ��I�!��J�Bj���BS�+S�a3K=L�!򤁢@Z�X�U�Z�KY�h{�$�f<!�DGx���E��Z>a���^2$!�D�7)z$ВB��^C���c�!!�dH.{m~=bi��9X1ah�t�!��ۻuQHcE%��<
�urm^�Q�!򤜾BY�5BB��+aJ����E�!�dE3�F%�æY�p��c�P�9�!�D�kQ^�srgQ�X�,�)��D�!�A�F�ӈ�6�Kx�C�I3nx��Jp�h����T��$�xC�� D/Dݳ�!VOͦ�9��_10E�C�I:Rb6�2�:��4��ڏ8<B䉅,��=�S��/ǌX�6�G�#��C�ɿx�T�2�� H����*j�C�ɪD
n@&�KJ�5{5OD�gs�C�ɐ�	3dƘP�(�P��)y4�C�I�kԩ8���c�����э-�C��r!+�K�lʤ����R�F}\C��	o���P��O�~�b�Є��{w�B�I�wRlu����=\
$ ��G2"�XC�I�,�6ap�d,�>�ഥ��? C��=, $쪤��I�"h�G^>M{�B�I�B�(��?[*���-PB�I u	(�k����F^�=��j�^{�B�I-�	�KW�Dxj�K�׸h� B�I�e��ܠ�H]V�N�	A� ,i>B�	�!r�t����bp^�S%F
�6�TC�ɞ;V�9� �5jbi*g��f��B�	�i�b,��Yz�x�K�;@�dB�ɻ\�H,ۂ�R�*��c�� �bB�	$ג`��BR���raO5��B䉯�*Mb�-�ri�Y�A��$>�C�ɫv>�5 G�V�6��-�`��~IdC�I(Y{T� Њu��o�2�xC�ɟJ��� �VA`5�Ҡ�0\bC�ɞ.��m�w��.���)E�X`�@C�I�c����tmV6x���#v�@C�	��R���'^ �q��a�hC�ɩ-$
=��͵s��B�$o�JC�	A�u��C�5n Kf3-aNC�)� �\�v��	Vv�0G"O5^^�#"O���C*IuAU��"_ ٣�"ONq�C"�`���y��	����"O�`	ՋۖN����e�m��m��"O���ÇS�����MdLh��"Of!�%įt� ��A�� d9�'Ĝ\@��
6⸳�MJn��Y�'��(xWeΦP6�x���[��*�'��X��G�i\Ĕ+����o�f0��'9���֋��b�٢�ԩe���'!p̩@K
�K$>�*���v�
���'�� 2�εU�v�'�y�0��'���"`G�[�(���qs��	�'��љ�m�=�F��v�m>����'�l�WoQ+h�t�H�臔c�`��'ڴh��G�g.X{e�������'�\�W�O;`�P���9{R�s�'ƌ��j�,��t��I�h����'�Uh�F��Z�&�z#b�!kQ(���'�M{� �� �>y+%B�5����
�'�\P�3��4>��2�.�4;�^��'v�I�3��
xlR�Ka���� �'��Y"��3r)0i���ru��'�� ��Ѷ\�Nu�˟�q���'�,\�uοK���� 
 ��Q��'¸k3a�kVz�J!�F� A4{�'�|��� �8#p�M���SM�t:f�B=*�qO��� ��?
��!M'�$��"O�`P�k'a�&� 6s �� �1�� 4v
�� ��7K�, �q��e�V9�cO���|�d=@<Ps��>c\�� fÿ{�
�:�O��PdjAEcaR�r)����S���Q��GB$HDx���  ���7u%�8�$��4_��i�R���Z�쁭�!��S�d�"ȉn��o$X��*+L:�{V�B�;�,�7ƃ{��������T�t��4V[쬳��� Aj�۵D�%��ȓ��]qsd��� =���$n����QJ[5A6�i
Q�jG�}�f����Aq3D3�Ď��U���ΤT����Fݦx��Qi�(�i��d�׉�P������ϧ�0`�P�2`�z��̑[��Y�
�� r<3f�a����/N�?�d�@U�L�t 
"`<�o\.&f��ᵄ6Iѓ�S-�p����df��N@ĳ��P�)8�4hA�1�~"�<��e��'�K��,b`��9
j|��n�=�Bp+!���,4�� &G3?�^�ۑ��7��>��f�Z
O�-Ai������V}���K��"9�!�$�*��-��Ȅ�M�}���B	�06M����1I�I� p�"�SlAS��0}b�����Z��$�:���'
��{eϗ\��d���9T�p�	&��z��E�$�"���0D~P�I��G�--Hd��o�D�(�REՐrf�m 6NMB��(ذaӝ�O4d��ʫ#��t��l��1���ᡏ��U�ࠫT������O���Gܧwǲ��~��L�v+��+!ސ���?�<�ǪN�m��<�b�(k����S���)i���� � }��H�`DI�blrgϯ�\�(�-�|�<�G��h�t�kgN�4�Ƞ#FE�ɶm 9�Q���b�+T��n?a#H�8`����h��O�S|��L�?/����M��I�bD$:r��e\�x0�J��^)i �"�~�b��
Q�X�}�OZ�#�/�3.��A	S��%d��I��O��1g�'Y��	�g���JivB�0ybU�U�ߑ��>�L�\4� ��.Ϣz���j�)<O�4�w�Ρ|���z�O���"�	F�����x0f��0"O �J��K+&�������Z4jB%�|�X
_8t U�j�O���+0'|�y;��$����'��	��V�x��N(�5��c�j�'Z2���>�s+U�x�����T�+g��21e�Yh<yЅ��_[�R� �GzP(vMȣ"Y��\"D���Q�i� =�'�G�'ֺ��TjοY9�y2��$Ѵ��*�}��	=.��Z��aG�\P�%�y���[K�[ CU>Q�x5S��Z���'�|%{�Z���?� 4m�DQ��8i��*6V� 9�"O�b��E�U�Ԉ�ĩ��JtVY���(�qO.���Y��;e�(���Q��
<zƴ��:�'b^�P��>�%OR����ꑔo��M�ACuH<��+�ɀe+W]T8R��P�R�Ƭ�n��p?aU���Q�鳆��*`���.�Q8��*�ڇA���BЛ�DB�G��?�4q�,TB.��'D��B�@>p��}z��՝+�6�g�/}ҀK�?]LE�wN�_�:U\e�^?Y���G�5�����+V�IR�&D�x�w��" ��+�"�EiX[tL%{��'�ڤx&��M���Y���2�y��V�%�b�����JTp�0���Pxb9�����ōA�2����G<rTr,�Kv�RФO��p��V�5�����d�/p޵���A	x����<	�x�&�* �5�[~~b.�>V��MQC�t���vFט���SEHX0l4�Q�ÜL�4�J>Ҙ��A;L*�Q�Ox�SiN�s�X0�L<a�R��$�h�'�$ �bGx��8#Ӯ	n\ZA"�'B�Y{�lL�.|�`�N2}D-�C�5���g�.�bI�i��8��u(�Do�����R����*1!ҥ"`($��b�$�>l�h�)樅�f���F�̋F.֟��I+'1����͝-��gy��G�pl�Jh��\lY��e�0��<A'(�]nO��z��M�KN�B�j��r�Z��ԫ\�%>������-�a|rc�lT��M�H��@@��p=�e��n>x'U�v0��t �F�p�a�G�#��A�吊͐x2	�Y�TP�Э��}��lF"��'ޠ1����%Vb]{�C	A�q��uB�FW/��E遯��b�>���"O�ht� ��oH�4��F�	�zĐ�α/���[#�i��#}�'��=�&@Z1Tg�A)`I�;1���"�'�f�!�ׯ�P�1� �0� t�N�v�Bq�p�[S�B�0<aD������;A���⃈>o�x���N#��p��]��� s�
��*�� X��T�&g֗L͢���'�Ш a�G[�8��Y=XXjP+OeQ���0f�nIɁ�92 N0�VGP�7K�c>�j��-�tK����q��+D��w��t���!E�N��J*F�x$=)�Șt]���I/V�l�� �o�R~�%ԇ_�3s�74�5+�gĜ�p?Gg��`�M�Z� � ElY�p�V�LF bԨ��MAVȎ�[�oă;�t��'4�B�J�Hz���՛[������D w����g�	ouD��5��I2�z��ضV�`s��L I����-ʭ8��ec�'I����";L���-�:���'�刡��;K$t��I�'����0�ю$b�>IaB�X�A~�tUc�]K|�`�e-D��*��3k<VHP�AQ]6��%�-0�T-��#E��x%��*'T��O��-X�x���<�L����Cn��s���p?q�T�e�T�Є���$�)��#7v��	�IK�V,9aB2J9����D�4>� ��U�͉eE�;:Q�|h �BWx�u�^\�S7�ԭ���҉�xd��K�dI�B�I'G*!J"BѼq�$Z���l��	�ꑫV�;g�$��h��41P�ߔ!0�Ͱ�+��:؎ȉ�"O��s%�Y�j��j�3�t�I *;}.�5e,���@4��$	�'�t�)���C�>Y!V��/8��n��&�xq�͔0"��\��)��<�P�̗7,�!�D�	t0n� ��{�H��g��M!��1H�I�EX�Aް� ��"F5!�˚>�`عCJAIa��D�-8!�D	�J�����2CJj�́. ?!�D��F9��)w��T؈��$.��/I!�$"xn�Ix�*g��g��OO!�˜L�P�Y���*����f�J5!�$��?VL���mDL�����eE�!�$��b�J��wEGsL����E�!�D�C��Li��9�(�S� ��+�!�dV�$�<��rA6#Έ�󥏠K+!�d�5W����o��D�v��ꊣZ!��l�F�0�U�o��e9�ˉ6�!�$\-�(!6��4B��%�#ʝ]!���v �4k�)��y�.�Zu+��.1!�� 4��e��H���z�
��֥H4"Ob�p!OR3Pj�02�ʉ�[�8S�"O��� ��r<�4(�,�*���"O���G�!h �S��`Ԯ486"O��y�bX�$S��J�Jϡk�Դ��"O�S�35�(J���!�����"O`!r���{�����%�	-yTɩ�"OJI��D|鲢��wv̼��"O�̙�`��?�P͹�		cp
�e"OfA	��ܛe�r�Ȑ��p��y$"OT��!k����H�+	?"�Е"O�)�燔$%���+$��xC"O� �'��l�-:ԋ.�"x��"O�U�B�<7��J�1��@҅"O�UP��T.�0��6&��ԁ�"Ob��dߗC�ͳ�/�F?8�zd"Ov�����Hб�nLp�0�"O�d�-`Nԝp����x�@�}�<����-k��Z�D ���r�
P�<1Uh\�A��DʷFK�M�i②�w�<��g�B���!�	@����t�Qm�<y�BP=D�����?V<a�Kw���#E�x
���=/�E[u��3U�xt���2D�D@b�O�~�vi����Tm`�'1D�cgH�|@z��!��3DR0�)D�$qs  �x�0��ͼ8{f��$D� j�b�< *2�9g� ;�,� �4D��9�L�	"8�Iw� ���F1\O� ��ԇ��,�d�`���bS@���A	'϶⟢}*��1I�N����I�V�]�e�2\� ����IJx�	ېn8\	�g x�2�סC!����C�@{С���M}��t��DC�g Ȁ�Wi�FfX3p �r�8ZF���d@(��0��V� BY�nY��b �'- �3�ɳ+�� ��:�j���hſA��(�,�S�b�$3Y]���h�0|���V�AK���OY)f�����<9��_.���B��n~����}a�u"@�*23b��rH"����WF\& X�s������|��I�g0��ԁ˓a�:i"�!H9�LH`1����L�"}a��F�.z+�t��!>M���4�bol��O��ۅ��$ �֒O1�ne��˜VAȽ�ր�%���{���[�48���nM�Y]��'UQ�4\>�e��^��3�Ę]���bJG Y������3GB6��0WD��Oq��7�)T�X���Y��'*� ���Q�lJ���Mߝ�M�e�?�j)�ӭ�|�7��-4�x����<`,@qjD"N80�b�
׸i�3���N4���O���Ո[?}�H%���١Jy�ش|�a���F�^!) M��O��>�enN�U� s�@��^�%��(��y��՗S��	����!'`b0�CC��y�#Hs�1����#r���y�b�x��庐eJ?5&��B��y�d��h p  ��   �  4  x  0  e)  �4  �?  K  QV  ma  �l  [x  0�  ��  ��  ��  ��  �  G�  ��  ��  �  \�  ��  S�  ��  d�  ��  b�  ��  � > � � � �" 7) 3 5< �B L �T �Y  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9��CZ���1.*��5���#D�������=9js����]>+-B�I�L,����ơT� *S"0G��B�I�<w<̉@���R��Xrȕ(Uv�B�	�n�t�hՈ7Cn���ӳ;�B�	x�Ψ3�E�V�B�ʑ�ޕ-bB�	�K��� L0B��h�'��O�`B�I~����b��L�5��£~�B�	�0�dq�  -Nz����� 9�0C�0>a1%
�y�N���.M7@B剖+($�w������Ο&|`!򤂰V�dS�D�
��PZv�I!��"���㰁L5=�����	�!�ӄA��a Q�&�ʀp`�0#&!�$\(�����N*�Z1�f��+%!�D�J�ݨ�H�UwP5hd�	!�$C0�d��#��1a��ɷ*���!�$J�gÔ�[��,;�2	:D��J�!�d�c�\���HOOj��q��o�!�R 5rZ@
T�� ]VH�RbY��!�dI�{g)#��MF�EQ�J�7_%!��= G4i�� �<+������5�!�D
�[�T��"D�*��Mr�N�2w!�$�aFڈ�&�ذM�t�D��l�!��.a��To��6�F|��,	�v�!�DQk�m�D"��W���wN@h�!�X��1R�/߽`v�S!/Ìk!���/uӦ&�(__�Ո!�ǖE1tܙ�I�X�Ļ��̓�!�ԉT���k�E[*E������6#�!�d�zr��h!ꖰg;l\��cT�t!���k~�X oF>@����c�#�!�8H�Lk��7�Fxk��R/�!��Z�^l2��^ a���Rf�L�,�!�$�� .!���"S$�*�.��2�!��0BYڨp� �:8P���KȝW�!�*@�X�Oފ?g��ॠ_�)�!�$�P��+D����z�� E�!��  �!�O�M ��#Y��"�8#"O<��"��5Jf<a�AmJ-�Xt	U"O0�8��+��k�삓���"O����HM6��JB1[��ЫD"O \�!�Ðq����g)B�6 ,AJ2�\x� PB�P*Ybk8t H�$D�� ���'-B�ր]�h�����.8D�t;���w��y���qa����+D�����$�!��J�q�Ġ��k+D�D3U��
u���9��U����y��;^t�X�WJ['�z�22�ۮ�y�o�+q!���d�$H"��y�I�n}['zR������y�A�?��pDkc8d����B3�yb�
�x�*�Y&�%��1��O:�y��\�`�x�b N�����+��yb��,h��i�JF��aVl���y�eɊ�lcP%M�:mtU0�E̾�yb�A�U�͑�&ǘDc�!iv��	�y�n²vl6�!�5�>PVaC��yEF� U����Q0CB]Z2�\�yr��`�й�Z/���-�\B�ɸ$�q+�����X��BDz�fB�Ix$!Ra�Л:q�Hx�D�-L�fC�Im�^@�a�D:p��ș3&"Z6PC�~�"�:'HIպ��1��0� C�	VQ�!�)ǝC��3���G�C�0e�y:p"B* P��D�*͸C䉶X�J	K�*�$v���	�k�'��C�I0�ȉ�c��*�"U	�h�
�'�} �A�5ΒA��V�-�1@�'>|��"�F1%
��	�-4����'�^Mir"�#*Wr�Ф��; ���' 諁nÄ�̂e���k�'�j@{�a�i����b��p�����'u꡺�i�K�IAa�D67���'�`5+`�P�{��c���B�F��	�'��E�ũ_#J���ȓ΂g�Q 
�')�	�2�؉kQ �E�q�pU�	�'@l��A���b�t.D�s	�' � ���ʹu���:�f��o�NYA�'�@Ц'�u�����M#_�����';j��s��z:�yZ���V:j��'jQ`u��(&�%; EKI���!�'�:��i��m&�� �Ci��B�'�Eڦi���
PӇG�7P:$!�'�<DaS#��x�E�K-Q�P};
�'��0#B[i��S��5����	�'��p5�Ëi�&���$�8oD�	�'�r8�,	G%��3�6��h	�'xڸ�@�Ir��+��U�<��`�'�����8M���k�(�3�\�	�'F��c
ցn��9ܹ!G�	
�'�F(�A`�Nn��NQfS	�'6,-�ѩ
),�p<`1a
.&�H��'�=��"��'�,a�탸(�L0�'j��1._("�ݺ�E����!�'��� �o��yp���F���'�nD��K5�
iʶB&-��}��'�`Y*��C!;�Ⅹ&
�nlx�'�,T�� |>�-JS�V��bu��'0�)m�\��}��a�/P����'����j�uM.�ׇE�<Y�5P�'�~��JI�Lx���;¨���� ��x�@�� � #� $h��'"O��B ��D�2�$I�r
�{�"O(�$E��jX��豉�4_���;�"O�zW#��3AB�a�H�o�����"O��#�i� oD2-S��:k�����'2�' ��'��'H��'��'�9)�Z�����F�
�+b\8�0�'!�'or�'�B�'�"�'h��'/6%0	�	d;��3�J�:���E�'�b�'H��'���'R�'���'�X�G(�g��!sc�Q=C�ybV�'���'mb�'���'��'I��'�ʑ9W.�����0d ����p��'�"�'}��'���'��'���'��Ԡ�.�Pق��2-K�Y���0F�'�B�'"�'�"�'���'���'������щB<�գ��-��*v�'���'�'`r�'t��'���'���´Ҿa�>P�pc�`�E�E�'�2�',��'s�'��'���'�`m���:����G�p�8�3�'Ur�'*��'d�'\r�'���'[�YEF�!G��٨��$d�$8�W�'{B�'��'���'���'���'u��a��_3Y�b��֣�1?�u�����I���I蟌��̟������۟��dCܮO*̽x�A1	�N��Bϔǟ���̟x�	�d�I��������	ş�Z��澱�$M�x,̰�r��ڟ��I��H�Iڟ��IʟH���Mc�Ӽs�O�����̉�M��eLL�a����������Ц�á ��{1�8si;����Jl���'�b6M4�	?��D�O0qk@c�+jXi�� >FqӤ�O���Z9��7*?Q�OU��) �z/b��CgAvqʐ����)��'p�V��D����%Ea��c�D܂ ʱ�CyL듣�d�Of�?�����;��y��b�����VlI��?1���y"^�b>M����͓��9`w�\3�dq$�_RY��y�l�O�y���4�t����W:0���V9 �(� G��<K>�B���O� @�/� @@М�&n�-[ϜA��,�	���$�OP��d�L�'����\�N���h=Z/��8�O0�dg�v���iP��?�*�O�y*�íP�v0p�A5���PI�<�)O���s�<r�I�TN�2�*��$}lY�Dg����ثOVʓVB�6�4��|���,.����J�"T���70OX���ON���=|q�6�'?Y�Oy���J�aj����{c������.;:�N>�(O1�1O~�
a�9P!�L3:�ި�t��8�O���?1����]:%K�-�Q,�^��\ѧ
�&��R؛-k��H%�b>9f�@�2���/��X}p��KL*��|y�E@�z�(�ɮs��'���.���C�Ȗ�W7y��Ǹg=�����M}R�'6�БR�v�R bUNG�!��傝'�"7�9�I!����ΦY
�4
��j�3�D`�#سy�<x@�Lr�� �i��O"�R������<���ֿc�̉'i��h�a��-W�V��W���<��,�<�� /&aڰ2È�����*O��D�^}ʟ\�m@��
1;Luk�
�A�̄�'Z�� K<�1�i��6=�B5AUg���bB�0�"A�02e!X�*ap��4$�\B��������5���t��yIG��D�����.��-;V"<�2Q�l��ϟ��IF���	u��L`V�� 6p���5���I}��'���|ʟ<�����*i�� DP�6������(+�0|�i�\(������F?L>1��O8 ���0��-�P�B<!b�ibVy��C8&@��zE��`�'R剦�MÎ��>��i�8��מ>rx9c�"U7Rrt`�RLa�2�n<*���l�r~ҩW�>l~%�6Rx�	3S��ac-ڛ�|�c�Q:Dؘ�	Wyb�'���'A��'��Z>�Vn��Sj9�!	! ��<�a%�����O �d�O����̦�:`��I���|�6:��D�XV����M���|���
��f���1�4�yR�_}v�5i$H�C��!�F.�y"�صV[���	�y�'_�	ޟ,��>l��e�`��CO�@���b�����џ���Οȕ'�ꓜ?����?�bD�.L��&ϛ�V4X1�S��'I��=/�m�r�&��Q��2.�zm�q�ʲ?�l,��fg����5m� ����m���'��$�R������'�R��fD]�%�н`B/�>�V��2�' ��'���'��>��I<	zNLj�O3�"���#�*����I���d�<�4�i��O�.�:��a�*�*�,d�d�ش��� ����LX�Kٝ9��Ԣ«-	��k<N�0:���e��&�8�'��'���'Vb�'���;�f��~d���'R�)�fX����O��D�O��$7�i�O.��/1,kN"��0V����]}r�'�2�|���LNv�V�P���!�v��ǆ8��5�ul	��D�k&"!K��r�O&˓\bD�zFm^�m`BqA����,����?9���?A��|Z,OҀ�'���2(]��*����+Կ�y¥r�@����O����Oh�D֪鈩2���.�]��$�e� !��l{�z�t�Y�*矒�>��=� ������a��Q�|P0x2D6O���O4���O����O2�?1�.�4q�B�@��|���џ��	���I�O�	�O|qm�_�I�PV�h�Ad�z\4�APME:��$���I۟擫A���m}~B#�#�l�� ��;VE�!��d3}����ݟ�cE�|�Y���Ɵ�����e��2H��p��-�2�t��"�ʟ|�IMy�m�>����?1����_�B��Y�V��P$y c�͓Ms�������O<�:�4������RD��x�
?$yH4! n��Z�f��Dd�Z�"�r��������BI�ɱ��e85)��]��98a�?qRI�	̟���ܟ��)�VyR(mӸ	z��O�0z"|�g�;(� ��C?O���OJ�o�@��c��	�*��t�t�Q`*��q��;4�]��L�	:g�(�o��<Y��M���@���1�'�n�(�(P8*�\�ٲ_�@^�	�'���D�I���I�����P��l�4l¸R�㚘*��#@`�u����?���?yN~�3:��w�6��p�;:���Ɋ�}۞ �u�'g"�|�O�2�'Ed�ˆ�i���ڨJ��U����4JH�\!����'ܪ�UnS۟ zW�|r^���̘�n'~x��d�.
�8�/�˟\�������FyR��>9��?���� M�g�� E�Z�Q�0�+�I6����D�O���;��Z3���3GΜ;P��W�Q&�ɜ9C{���F�b>5s��'L�T�I�|���Q��^�ROH)E$	#u��I֟���ܟP�Ix�O��m] u�v��6D�H9ְC�m��h�>����?���i��O󮉟"�&�8��-�&���h�9��d̦��4��f�"]h�&:Oz�$��
�I�?=a�K1n�=��f9��13S���c��'�������ן����4���W�@1b���$39�|�%&UwV��'�\ꓶ?md��d3�)�O�%X�`C#��d�QՇE �z�By��'��|�'����R��Ag)<�^X8�F���`���"
tB)�+OX�;�c��?Y�,/�ĸ<yj�����7Yz$,[֮�&�?a���?���?�'��$�L}��'�J�B�@�%Y-�T"!�	�b�H̘�'g�6�$�I��DPӦ�+��M���·H(PːlE�9�<iJd�E1&�a�t�G�0 ����<P�H~���ʠIAbm_�Y���1�	v:L$ϓ�?���?!���?	����O��!Jwg��te03��Q�X��'q��'�h��|���1���|rѹ+��V��?�]A*P�U�O���O�FS�Rݛ��T@�- p�T��F낵e�T;%iA��"=��'�.|'�(�'�"�'���'���p�����IE.�*z�xq�'�bP�`��OT˓�?�(�,��#��X�м�5�#8�ڑ��(p�O���n��%��'>A�<�R+H�i���.X�rK(��͓4��ԁ��*��4��P���k�6�O�H�h�~���:��۠! }�ת�O����O����O1��˓Z�&A	YhLujZ8[�
�S�FZ�y��'�2�p���D+�O�!m�R�T�%E�e�4�����(G�h���M��L:�M�O������3���l�<	� ݱ	�@�僟	��]��m��<�(O$���O�$�O����O��'��5(�DW�Vzqz�[�HS&]�\���	�h�IL��̓����1�);��X)�d�	�3ae_:.�fa�O�O1����Ѫa��IQ;��;��Û��v�ۥ`�@%�'�Ι� �D��t
V�|RV�P�Iџ,��ޢ�lZEk�4:T�v��ʟ��	���	}yn�>���?	�C�P��;|=��y�+{R���I�>��i�x��7��[�UE��Z��U-4�-�&���^H���ZR,�� �W�LX'?���'�L|��/by�taf�9c� ���ʘ"��	ڟ��Iϟ���b�O��@�%��Q�qOY�'X!� *��j}B�'��fcӼ��]6$��$B��)j5���&�I⟜�Iџ��tK���'D2T��&�?mB���1ň�g�6C>|����&k�'A�i>Q��ԟ@�	���	</�z�Ye@�=����ƣ'���'0d��?!���?�K~��Da#��F�~(I� ��7
���Z�<��ݟ�%�b>i��c�Ƚз��.`N\�/��q����O1?�Y E��$�"����Z�Jv�`�qF/z:��n�"yڈ��O
���Ol�4���'������X�a��;L�7���=��Y�d�͟б�4��'�ꓡ?A���?1Fh�SE�Z��Y=�8�!`�5���Bܴ�y��'j�9����?I�O������&B˨J�1�D� K�ʥ+G;O����O���Ot�$�O��?]p �E�fI@��
$l#|�e�Dy��'� �S�'uӤ�OH��4cT�0h�]��]>(EԈ�e�$���O��4���x �z�`����X��G��v�Y�+�vl`�2yt��`��y2�'�2�'��	C�E>:-xX+1xY� ��\�B�'��,��$�O����O�˧d	*�kH�3Cޝ�O��+4A�'�꓋?i����S�T�Q%�P��uN
��P1�M�GtU#�@�[֛V�<ͧ�8�Ij��=6b�9(A�(dɒ�ᇀ��PF���͟���ş8�)�KyR�d�8���L$K#*}��A�;3p^`4O����O�oZJ�7��	���z`k�~Y|�p�M�	��@��-E�����*�TlA~"�__&�`�f�� X�"v��J��%�"�	f���!2Oʓ�?��?Y���?����)�֘h�\���+�e��ifq�'���''����'I�7=���
tA�8�� �)Cwʭ����OP��/�4�~�d�O�P���z��4�Xd��O��A ΍�	�^�	�~�L���'���$�H���4�'��m&	i0�`�  ��-B��'��'�X�0��O"�$�ON���-F>h#�)$.��͑5��#���0r�O��$�O��O�X��#��L���Rdi/u(�H3Ė������$��m� ��'I��Iߟ�O�f�؉��� bs�D��P��͟��	���F�D�'��䋠)�1> >��Cg�^���$�'�2듸?��fI���4�}�R�E1W�,�5�Ձ"e� 0a1O^�D�O��I�*�7me�X����LI ҟ�ؑ��d]��� LX-U��q /�d�<���?Y���?!���?A!(D�P�ɍ�E�1a� ÷���t}��'"�'/�O��+}5�,ڡ%N�R�8ŅM�n8~��?����S�'@��[���5>*NiAp�=a�M�� ū�M�EW�K�l�,��/���<i0¥g3d���.�4���g��$�?���?Y��?�'��$U}��'X^���g�iG,�E+�)��Қ'�6�)�	�����OP��O���CS(D�>t�3A��@�2KM�oZ7m9?Y�"̬=���I0���1�1�J^ct����5���j��h�0����`������@y�����@8��a!ą�^t��ba�A����'NBö>ͧ�?�i6�'����P�B!,�2!"���:�B�{!�|��'+�Ow����i���:2�*ă�"��0����G&�c�ra��e��8("^�y�OS��'��%N�B��=["��u�~��K��&iR�'��I>��$�O���Oz�'4:q�� 
��y�0-P�X	�U�'vF듨?A�'Љ��I�2U�tr�-��J�u����7�2H����"�"
����|��b�O<K>9ЂIh����ìα$�A2���?��?q���?�|�(O��mZi%Ri����4C��T�&�ן�	��M3�b�>��:���nǛy��G�U5S}�q�'��B;k؛���py�M>x��T��ky�|L�e�7g��(+�ʴ5h�����O����O��O����|R�F���X���V�~��Ԫf$tS�Ioy��'��nmz��pO�.L�e���9�JIS����M+ŵi[8O1��$A�loӴ�ɂ_
i[F�R�LqpV��!KT扷e�m9��' ��%�h�'r�'e����ʲ$��D�"&Ԝ�C�'�R�'�BQ���O�d�O��$�g�� �AE�p(�iVB�	|r� ;�O��D�O,�O5�"D��b���F�~H)`�>O.���<h�TB� v��'����[?a���H�DDФ1����	��a��?a��?���h��d̝*ۦI��L��Qe��y%��*Fb����F}��'��n�"��s�h�0B�2���D���oy��	�0�Iٟz��ɦi�'d0����[_Z�IQ:�B���ݏ
�� (A�9����d�O���O��d�O��ă ��h
c�ϰ";�UI��J?���Iҟ,��۟�%?!�I�(r �ҋ�J�l�z�$�<��]r�O�\nڼ�?qI<�|�!��'�Hpz��D���� �/XD�i����d_$P�l��O��C�ĉFjH5T��},p�q1!X��?y���?Q���?�'��z}"�'9
yI5��2 �@��*(�:Z�'��6� �	����˦�����MCq�Z��č�g��n��g�˗	��� ٴ�y��'ӌU�C��?��_�\�S���Sf5aP�j���=t���nn��������	۟��	ڟ��*���c��ͻ���[_Y����?��?�wQ��'�Z6�>�$G�y��("�͊Z��a qD�J�r�$�d��Ο�IL/P�\6M<?ّ"ٮY�Z�@+�3�@|	 �@!����u��OF�xK>�-O����O����O�����3���ु#	_j�����O����<-��Iܟd������OT���N�R���g�+*'*�x�O`D�'G.6����%��'%S<7#Ő)2L(J��B�x�� r2�!H�P� #���4�a:��ГOj�q���{�0�v�O#��R�e�O����O2���O1�Tʓ{<�ΜF�V�ñ
��� IP��yBZ��ڴ��'���P�f��*=U�AW��9���gE�DgL6-��m�O�զ]��?��:f*.��_>��L1<(�gR�,\���Ŏ�+}�<Q���?���?	���?q+�Rp���d=�D��3^?H)b�ge}��'��'*�Oblq��nXDm�9jE*�O.ܡ���cF�D�OV�O���O��T�orj7�a���7�؆I�漊af��"�I�oi�h�m�.b�$/�d�<���?	�� ��� J�2蚬�à�5�?�����ߟ�'X���?1��?����}��c�`�x��� ����'���?a���|�2Ռ�����3a�0ϓ�?��@V����3ܴW/���?�P'�OL�d���*���拏,`jaL[�@�D���O����O��d!�'�?��ӈ��*GS�+"��ځ ��?��]�H�'��7m/�i����S�dt��"IDOŘ�r��e����ޟL�I�Y�mZ|~"�S!f��=�g�? ��م.ݞ:g@����:U�l9�W�;���<���?����?��?Y�ՏI�  ��ƊA��13A���NF}"�'=��'2�O>��ٽF�L8ꠣH�窩U
ȣy���mD�v��O�O1�,�*���$	���fD�e.x)����"N�L�H�<��D:~��DB�����D��|P���U%��
��H�!F|�$�O��d�O��4��ʓ@���˟���*P]}�͚^#0�]*�JV��cw�d�tѭO����O\�ğ���ɸ�+�b,dL��M��P�w��=O�$D�"��M��O!�	�?��]*,��M�Xh5�u�[5�T�#=O��$�O����O$�$�O�?����U*�����Z�g�J��"���<��ٟl8�O^��v�|"���N��i�cåM�:x�$�ӘZ��'�r�'��ؐvs�V?O�dX-��PZ����rBֹ ��Įj��cǊN��~"�|RW����̟��	؟|���)q�6��B� �m�'F�����Qy���>���?a���Ձj�p�!3�z���K��I�����O��D'��?��?3��BV'�R�d4c�.M P��IYG�
��}�+O�:�~җ|�` `��lH�fG7��x���3W��'5�'��TY� Y޴!�Tɋw ύ2��5��F jT,͓�?1��]ɛ&�$ry�i�)��ͭY_z��p
M1AW|�����O�6��t�7�=?q���,#���I�����(z�4|����[�� �!��$�<9��?���?��?y,��)�LG.��XSw*�'�0��oB}��'�B�'���yҡa���Wc��:�H�i��I���[�l�йmZ��?�J<�'�"��y"���4�y2��y0���.:]4ͣ�a�7�y���.y"��	?J�'x�	ğT���s|�qFR�Z��ܡ̈́�>@4A�	֟l�IП|�'��?���?���ʤy�dfcH�/���$NC!��'����?����$�����^.!�(��ԋ���'C`Q9uƆW��(����~��'�(=��:*xF�i�� �*�P�'h��'�"�'��>]�I6:L9��K1tu�߻C� I����$�O��dW˦1�?�;=j^X7�n�Z9�v"��f�Γ�?Q�x&�Viۇ7��?Ox�d��iF�����V)ytI�&�<��C�6N^����@4�D�<��?Y��?9���?ل� w�X`S��)J��q� A���Ip}��'�R�' �O���X�K���)�ĉ�<����ӕt����?��'����O+��ش��0.�RM68P���.�3u:p�Q�Hy�c�8I���E��yy���!�-����A������'���'��O��
����O���c��M�L	��N#����+�Om�k��v@���M�2�'��%W�Eٴ��&�"��x �/�)h00f�i��$�O�16�����M�<A������`^�hMx)�ڏ
8�L�GA�<���?����?����?��T��	Y�P�����j����L��'��>�'�?��i��'c�L�w��?d�MP�02�䡉4&-���%�ߴ��S�#�M#�'�M�|�4����5N������(1ZP8��-C�t�d�|�]���	������pq��D�|x� �\�B�T)q�Gٟ���Ay��>i���?����F$)+`](fB@=�t4B��
+�	���ʦՂ�4Y����D*BJa�C"ޟ �����*��R&B��$Č�Na@�!���<�'=M4�$����I$D�񓪅��1`AE%f���y���?9��?��Ş��ۦq3!�9J�������F;,��`m���',7�%�������O�Qy ��XLx�A�/�&e���HT&�O�D����6�}�t�I-t���(��O��E���pҦP�u�L� 	��z�����O.���O����O �ħ|�o���|����@F����6��	̟��՟%?�	��Mϻ=ǒ�C���jI'HJ��&L���?�N>�|�h��M�'N"�����"~@���$�	Ϣ�8�'���⧤�Ο�`�|�T��՟���E�L�����\_xkei�����I��P��|y�"�>�*O����o��,ѐR�#�9a�J�� >8� �,O���O�O���ת��@(8@��L�b��3O4�D
�������(_Q���J+�OhE���U�� ��y��$3Ѐ�70�X����?q��?����h�R��4'��h �(C��������9:���T}��'B/z�\�� w,��P�\�4�@K�;Y@�I��M+#�'꛶@\�-W�����P�C��[O����rq*t�a�*�"#b�5��5$��'��'�b�'+��'{�X)�@ͦT.��[o��M����V���O����O��$���Ot|�r�4i��c��Y�fc�x���gyR�'8�|J~
u�.`y��s'��s���`\�N	��'�#��d�DLn�j��m�ޓOd˓X��h3Bݾ``��91�m��8��?����?y��|�)Ofl�'������r4o_ vd����e��!H�'j���h��OHo�?)ߴ\�n�1�ʡ���c"%��1v�0PQ��MK�O:��c֠��r�&�����|p�S)wY:�Pƈ�
o�EJ$<O<�$�OV�$�O��D�Ot�?�s�+:Q����+�a| �8����������Y�O�ӧ�MSK>�%�\:������dD��f��-~Q�'Er�2�N�MC�O�A�� ހ��N�Ox�Mc�G�O�T��̸�?���9���<q��?y���?�����rc�԰90ΩC��&�?����D	`}b�'(��'�Ӭ�~qPP�57�|�[E(�s�`�Zo���M���'���IQ	=��0����$�o�&"���w�H>��HJ��<ͧ/l��Ą.�� ������\9g��h��3��O՟8���t���b>��'B�7��8�� ���#�NM3хX����O��ę���?a5]���4�l�9�C}��1���T�͞`�6�'-�6ǈ�B��v���hQ)�8\���*OOy��A�)JQ�f��m���٣IŤ�y�T�H�	����	��	埰�Ow�Q0F�K�"�⠃�#޺A)>�WC�>���?)�����<Y��ywσ�d�D�f�����)&hw>6m�Ȧ�iM<�|���� �M�',B��k�*#��%Q�H���"�)�'���0rk�ӟX`�|2[����ڟ�a�g��F���G�/�Re�o\ӟp�Iğ��IJy⥯>���?	��
���s,��t�\��`��#H�<�"Ͽ<1��M�@�x�R���x�Ff�)@A����L���:�^�s�g8����j�K��:���dz�ӉB�%��P;�%��#a�h@��O��$�O�D�O�}�;XwJi�g�2I�Nt��%ǕJ�~0��]N��vy"�n�`���% �����0H9 �3��������Dn�<�?9���'��#���?�;"hܒ-����g�h�@�sQ�'U��'��	⟰��՟��	͟t�	6#������ɽڠ�3�E?Z�p�'����?����?���df�}���ӢÐ�P=����=4��?�����Ş@�$���S=a��iNK�j�ؠX�O��M�!W�P+���~>�d/��<9���1���aN��k�k��?����?	��?�'��do}"�'�����1"���g@�[��z�'ђ7m$��,����O��4�.U)���u_�m��M �u�t�$�\=�7-&?I�)��ATB�z����7J� ��;怙1K+%��g���ퟘ��Ɵ��	����ʃSI
U #"O)P������?9��?9]�����4��B�Pmz5'���8�Hc/܁���9L>I���?�'[8�)۴���P)t�d��W�(z����{̩e��~B�|bZ��������I���"p�V4{3��-�? ���z�����(��~y��>q���?������X�6�p'��&�=3"I��<�ɦ��D�ঝ�����S�d�͞U�ƀ��`�/Ud4a�� T�YU�ǋp�	��U�擒%�$U�	>��9���-cQ\	CLW�`��=�	ҟ���۟(�)�Uy��fӈt��
20 �"��U"0�(��D�O��$�-�?WY���޴-h����8*oN}*��_ n���ۡ�'���M�bg�������O�6��T/uy�KG�eS�=�HԼ}w0��yrU���I �IП��	؟��O3�yHP���sp���%߫[ �g�>���?�����<٣��y���"�b�ӓ�W�@TP�XUD�$v_�7�̦-�M<�'�*��;�E3�4�y�Y?$޶� =]䠸T䒦�y�mۗk6L�I�KN�'��ӟt�I.4�pehӢ	|�H���b��%�Iߟ��	ğ䔧�\�H�	Ο�I�w�����O�2M���M�)����? U����4*d�Fo0��V�fJ�R���-b�P� ��O���>>�ĨCf�ɺ���&?�[�'������&\d\���B�� ���Z>Wʎ��ߟ��������{�O��é!Ķ�+Ѧ��dk
�9FE�.%h�>I+O�dl�a�Ӽ�s�kj>�`$�M-s�$��+�<���i��7�Cܦ} ��ŦA��@-Y�_��χ8x����G�Tu�䱷�֝a��'���'���'���'_��'��M����R�h�h�C�T}vA:�[���O����ON��7�9O��`���7�x�'�m;�X��'�L6-�ԦQCK<�|���
06?l�[dCיy�~��e
�{{`�S�c���D�)U<���[��O��Z�,u:��M8gtQ��L�6�&����?A��?Q��|�*O�'�R)Q�D+��BC��
\���Ѱx�R�y�⟜x�Ox�$�O&��ڮ��`��\�W�f�FPEUs�m��U���?�'?]�];����VE�(�:����)ft�Iɟ�����x��ş���f�'c��Xa-�=p����M3u��q���?a�>��i>-����M�K>Y��	�� b��?~�FaA�吂���?A��|Z��ހ�M��OT����-8�zD)Cm�dUʝ�a��R��բ�'�'���Ɵ(�����[����G�@��@,x�ݘp�'��X���OP�$�O���|B�ʋ.~��Uj7�Uy�.���W[~�H�<	���M�W�|*�|�rp�W-G��!ʹ;�؁�D�/J���pO��0����|�"�O�8�J>yuB�=��acfY"FW|�q(���?	��?���?�|
-O�=l�s%䐫��O4��MA:cIz�yy�g`���|�Oh�o��	
��cqcK5ռ}��HG�P��ԑشb.�V���I
ET���O�h�e�	�z��<)#����P�86u�d���<�(O��D�O����O`�D�O�˧*��ʖ�޵&�zE%��5S��� ]�<�I� ��U�s������c0i����uFm�Qp�����C���ӀY'�b>E�jX���S�? ���^=�NT ��Z!+$l��6O��#uJ���?�r #�$�<���?�s�ܿb���Cb���K�G�?��?�����Tk}B�'aR�'��Cwf�7q�(�AՌ��z�B	zr�dh}r.fӸX��A≰�:q�[)^�m�$n�\7��P�2<�@�5x�p�PN~��On��+6�Hg�֯o�@,jc�E4
(����?���?����h����(rͤ�˴*��[z���FIdk��Di}��'H�jt� ��Z�(�3�_�D� ��cIu��扚�M��i�7M��_QF6�e�T���k ��H��OP�h��Զ]��`�U K#)���3�+�t�	by"�'���'���'�R�6nt��+<�
<@6e�)�剀���<������?9ӥ�c��u�3�ԛ�LI�Bj��\���|̓���|B���!�F����2E�&J
� !�"��Ux�H"�7��Ę��`X���2�N�OjʓT����#���8Ą(�$��g�h�(��?����?y��|�*O& �'���N#,��x��!ɘ�ޜ2�ɀ��y�Ho�8⟰۫O�mڮ�?��4#����6؇v�\C�@�+�z�8��� �M��O�h:D�I �R��<����d�����#�Za �,�H/zY��8O��D�O*�D�O��d�O"�?Y����K���2ց��"dY�F�ԟ��	韌 �O���O�oI�I�q�>��� �=� M��-D��%�L�����Ӫ��o�~�g��0�K`�%s�H��
A�f<�*�)|?qM>�,O^���O^�$�O0(��� ��}�6��Zj=��"�OZ�D�<�wT���	�$�Il�4���e��&rl0��ŋ����V}­l�Fpm����S�t���}A4x�4S'Q�|�+Ӹ���"�%{0ab�X��SU�҉�a�I �P�Ä�+\.����T�F��	�X�	����)�gy2jӺ�;�$�+kF��&�ǀP��с;O�ʓ(���d�@}�|�j�`R'��J�$-ψ=��%���Ȧ�QݴvP�Z�4��䏪_�v��'?���us����5�*P�rFϯ�N ͓����O<�d�O��D�O����|��DΌq���r�ڱתQ�oO��ԟ��	��%?牿�M�;B�$U�� o<c!gZ$8�Q �i 6��E�i>u���|��d����͓
��B`�1a���&#�&!3v��)���OxiJJ>�.O���O��(a�Ͼ���J1�Ϟ�@@+��Od���Ob��<�3[���Iş��ɈD�\| a�G/���p��8;�F��?	tW�|	ٴ6=x��G�;��	Ic��"Pd���>���T3X����2y(j���I�|(x���?oJp2r�!;�d�i2�N�a	��d�OF���O��$-��3 %ͻ���.%V��Ŵ.��)�I���į<!�iS�O�3��hHC$B�6	G!3�����@n���M�⢛��M+�O�<��cS�����q �$�EKQ�Jݺ �Fa> �j�O���?A��?����?���t���/� NRx��C��`�/O��'2�'.��'^�IZB��2Lmp�� �1�Ȍ�ţ�>i��?�L>ͧ�?��P2�ч�
<wN	�G�@-b����T�\&�M�d^���c�:�������%#�b�@�ϙ�����'�4}����O��O��4���}	����<@tFߏ7]�̡gmP�X��x#��m�Dq۴��'3���?����?�4f�B���P"H�t�r��b�B�f2M��4��D��+]�9�O�O��-�8�H��*�q�P(9�y��'Mr�'���'����^>-��#&I��:��vA�l�����O���Ix}�O��wӚ�O���]8D�BCI�	8u��<wI�Ot�l��?���aK�ho�~~�$�?0gN�h�i�Y.�}�#�26��	��B̟0�u�|�W���	���	ӟ$�1�I�#��BA� ΚP ������I{yb��>Y���?����iW��b���K�EN�x{4d�(��	���dIΦm�����S�ą">9��c7��/f��@bogXX �#c��}z����V��9��Y�I�w��d����H��<��i��z)�	��p�Iן�)�Gy��t�NHj�O2�� l,-���;O��D�O��n�a���ɑ�M�c"U"^rX�m � Ր	R3ݨ'�i�"�ٶ�i����/,e���O���'�� ��qBT��4�Н�ß'�����ퟴ�IٟL�	M���Pk�j�O�W�ΩZ��Sܞ��?����?����s����D:4��F�6�B�@&&I�D�Od�O1��i��#g�N�	_�<E�5I(�<��,AG}��	$a�����OؒO�˓�?���S�l�Y�%;H6<�0M��&�1��?����?�+O�A�'���'��A.GV��vL((f4�r-[/*�Ofa�'�r�'n�'�v@�0� D�:�@$f�����O�̑uF޵A�.��Q�)���?�QC�OVR�L�(h���݀{��РEa�O.���OT��Oܢ}B��7��y�D�ԯ%����lT8h}\A��o���vy�@qӼ��]��e���<��P'^�6Z��I��M��id*6m��a� 6�=?S�]�yn���_��
u����O��$[�/��5<�UH>q-O���O����OX��O*tC#+���A�P�%U��S�-�<ɅU���ԟH���s���7l�E��d�pʔD.�iA�Z3��$�ƦiI����Ş'Vrh� 
�� �h�j�s�#	����n=	^�ʓyPL���O0x�J>1(OP!�$̘#z�0ѧ�S !ҶY���O.���Op�D�O�ɨ<ї\���I%[��,��^81J\��B��|]���M[���>iѿi8X��v�>�դY(0Z�m(�����D�C*� qd7�&?I��
�v�I���'���%��x-J%Æ2q�RK��
�<����?����?1��?����)V�V#�٩&��X���ui�'�r�'�2˨>�O�X7�6��1��ke���rA����I�B�Or���O�#{��6�9?q��QǢ�0`�\���C��O*h��e����$�ܖ'-��'�R�'om"��þb�sd��%'�4��W�'k�]�(��O����O4���|��NBB�ĩh�Ɉ� �}~���>���?�L>�O妵��e�u�|�a�@���FnZ�y���Եi�2��|Z'ȭ�@$�P;�O��"\6T8e�N�o6��� ��L��ӟL����b>͔'��7�?)���p�J5���aUf�H��Ŀ<��iO�O���'� ŋ'D<�� 0G"��RҪT	���'��i$����� @�O��5[޸��oX!Ը���&t:$̓���O��d�O�D�O����|� �W-�l����a��} �
փ,��������`$?牸�MϻdZd�#�I����c�[��xdJ��i$���3��I]>7�~���7@̾@��e�壐�."���'v��4�})���\�O�˓�?��S�(��'dT�5�&��ש
 �-s��?��?�*OD)�'���'�"�Cn�><�!=�6�9�%�(@�Ox@�'U<6-J��d$�h����Q�@��(Z�,��s�>?!���:q���&��'�$�䚦�?�q��2W�V�`@n�2�,�o��?9��?����?���	�O��?"���kM�2%������O4��'o��'H6M2�i�%ҡ)�� ���XE ��5�2l�6�a���41���i3�!�°i����4'2���O��Y(�:�r��	�N�XiB��G�IBy��'!�'.b�'9rBUzA^Q��i�"����c��?q�I���D�O��D�O6���$�x���uC�`��ݸG�'@��4�'z�6Y͟x&�b>U�C"#i���Lƿ_y$�iÌ�^��80b��my§Vra�I��'�I*�)k��
E�z��HK֚���������4�i>)�'����?q��D�t�ʄ���Nڅ�ʂ�<4�i��O�	�']�6��0lZ=�ֽYa��6gԂ�I׬ڡDW�1҅�����'�}��n�?��0��d�w@Y�)X�� ���5tw�3�'��'�b�']�'��֥�T�z���˓I� �Q�O ���O�9�'��7�M�N>a5AШy	VŪ�ԓ>�X�'��"V�'�x6�؟�I�8$�:6-$?A5A�("x��g�T!��H��B.4������O 0	M>�*O@��O����O�Ŭ�[���y�/ً?�̊q�̡�?����d�[}"�'�B�'9��I H N�<)�V��5II� ͪ�HS�I�M#�'B����W&{7�]����6m)��9�ve�sc� �|-�Qg�<�' ���F��;��J��L�;�6yU�7�� ��?	��?��S�'��F�=�S(Uh�n�S'���i���S@�p���'̤7-?�������O���@�G���6��fm�	��O�dҫ>�7m ?I�d�q���8��'�^ЪTr��D6�����k��y"]�������������埘�O�x	�f���uNv� �e
�*��C���>-�M���?�M~��$ޛ�w�l(���Q�q���0���'�Ґ|��$�Y�62��9O ��&���N��%kf�P3C)"�q 4O(�JE�x#�(D��qy�O��Dّ$Ȳ�0F@��}N\1��Q�Q��'��'�	���d�O(���O:U(r�
`���r!�H�&�3��-����O��$7��I�`��b�<CR���\i��>y���F��b>��U�'�d��0j�l!8��H�7J�*�l\VA8��	ʟ��I���x�O�R�	�+f�&$.}!D`��,�4f�>��?��ii�O�"Q��u���;$간���Ǎd�D�O���Oy`&fӀ�(!��a���P�RU�?�$�����\�RMB�����4��$�O�D�O&�
8s�UQe�0G� �v��/f��ʓ���ߟ�������J�(Z�9�����D�X�K�=A��B�O��$�O��O1�v�ఁȪ�fm��^3/%�����B�g����@��0	Âh�r��l�F~¦ù�T$��G�>'������?����?����?ͧ��$w}�'D6���+�%���)��ee�CT�'�P7 �	���d�O����O�i���
�����`���U�H�.D�7M:?YW��#`p�I �S��)+WaJ.�ZM�s�?J��3t�p���Iٟt����������r��T&�L�b O��:��RH��?Q��?\�8�'26�,����:\RS��С~�AVJ�
e]�O�D�O��ɡX*6M9?10.�]PJ��#��1t�x���Q��5�%�O�#H>�-O�	�O �d�O�B��I0RJ�� Ʌ�'�� �u�O����<Y�X���������[�T��fB���,n a���ދ��$�m}��'��|ʟ� LY��e�T���Ĝ	�B-CR�Y�Y��DR�~O�i>���'���$�4ɠ&S�*i!�Ȁ�����dݟ���؟|�I�b>�'�6���z\���Z�rU��8ʰ2��<�iQ�O���'��ȗ��x�!r&d�fᐪj��'�ܐ�G�i��I�D�9� �O0�'h���gE ���Y�i��	  ϓ��D�O����Ob�d�OL�Ħ|R`bH�Y�F� 0&Z�A�Nu@!�,$n�	����ȟ8$?牒�M�;o]�h[p�V�Z�1A�,ߍ f�l���i��+��)ր(-�7�~���ß!e��[�.�Q�̪f
s�b�n_:�⥉n�zy��'
�����Q��C�;]�}�ƃ�;F�2�'��'�I0����O4���O�3���0�f��GԠ<,{��,�	���ŦM�����oV����(3�VɹB���u�'bP���kʳ�\��e���
🬛��'JZ�F���Uv��H�9����a�'���'���'m�>=�ɅIN b� �$)�~��%���[rp�I3����O�����)�?�;�����$��'D�x1�cϐx������?9��M�����M��O��7�)��h t��(
#��3gB#tܒO�ʓ�?a��?����?�7��  �r&H=Z��G�y��h*OL��'���'R����'�6�H�,>̒��`Z��D�vN�>a��iz�*��)B<p�j��]�i�^-��@A�� R��U+1���h�ZҨ�O��zO>A*O��#���Al�yi�aJ6���K��O���O>���O��<�Y���I�a����b.	&j���P7۶�	7�M#��+�<���?	޴����c�^X`B�2@��`s�!U��M��O�"��A�"�G"���H�%HxH#��>pNp��2<O����O����O��D�O@�?�4��̚�����d��d�ϟ��	̟���Opʓ,1���|��5 ��ٳh��g�f<jQbڻQ��O��lZ1�?�a�LlZh~R�� ��S#�[�l@=�e�[!l�X�4���8�Q�|rY���	����I����#%0�{�!ؔUX��J����	ayR/�>q-O����|��$G� �\���
	.ڌụ+�<Q��d����4m��S�D-�8(JG䙲?�ԕ�v�Б0�P�ӒkȠLݞ=�@Y���( ��,�g�I�3����,�A��P��lX�'qJX��ȟ$����D�)�myr�eӴ��#�Ҙ[�*y��\�"_Px�R8O(���Op!l�J�	埬K�O��l�8 t�̻�DY�:zDk��G?�	شx՛�`��/K���ԫFM�(;����}yR�̏ƈ�*��I�������yr\���ϟ��������ɟx�OĬ�zr�� ~i��9P�cz��K`ȳ>a��?���䧧?IQ��yǏ�;���{ Nz"�mX2FK�"�'�ɧ�O�����i��N|��@efC������<m��Dtf��'�'�IǟH�I�5C�UZ����\�\����I.Ij����|��П��'������O0���'ԯ�Еb7J�".@,���G3�$�O���'�|7�-CL<��C�MY𤒦��)LTQ���A~bMկSQ*e�1��
5��ON,y��5�2��^L8I�	 �J����IN�[G��'��'�b�؟�$�X*(�2�A�C�&w�M�sfJ�èO ���O$en�z��՟�_Rf���j@��3��2�z���������0Ae'�;?q�g��o��S�#~�@s G;@�r����6�Q'���'�2�'��'�b�'8P��e �
$� ��įOb3�!�W��C�Ol�D�O��7���O�xB�� �l��U�fL-�F��R��g}�'�|��d�Y�{�0����"Th��I7O4:�@Q�i9�˓=O:y"�!���'���'��R�
�5��rYC�6i��OBɟ ������	���Cy���>�i�
����G�~ ։ t���g2Έ��@+���|2�'�T�p6��jfӢ�o*��34�L������st�D"�ܦ%�'{�}�akG�?�:�����w��QrH�@��!��L�8�˙'�R�'[�'���'M���4DW�!Ж�j ԱI��<�L�Ox��O�=֧���'�h7M<�D�O���]�&�J���iUB�e≝�M;���p!�6�M��O�Qj�nR*X���ШG+��3�m"F�����h�O˓�?���?���Q��蓭ѭu~���l
��OB�ĵ<�$T�����(��w����p�>�;D�ːq֜�h� ���W}*p�@=�IG�)
q��8�p�i�Ȗ#J�xU��AJ���@�D�V�r��,O�iQ��?��2��	�F�TZToͥ8�p�i���{.�d�Of���OF��<i �ivN�iQ���x�\X�CV�h4���'��'Yf7�&�����F�3��j[:l�nؓ��)Ŧ� �?�޴.�@<k�4��ݵi�1��w��T� |"��>�ʬ�BE��ϓ��$�O����O0��O��$�|��A3q��h���Ш	���  ǵ���ݟ@�	Ɵ�%?�I��Mϻc.��G�yj�	Bč�y�`;��iX��-����3Uz7�v��G	�~�'hR5R~vx�y��@���x�g�E��Gyb�'�2�ܩGLZ�[��p� ``Q��%���'�'��I�����O���O\�����	 hJ�B
C%�����%�����ɦ�����S�? L�C�&�@��Q �P�yy��:�����T(��;���k�Ӆ'r��� �5� n��5p1�U�)J�0��C��	՟���؟F�4�'q��S-�V.�uڇ ]&>,����'����?q��	֛6�4��d��ߩU��������FL�������ߟ�oZ ^�o�Q~�%\�A
H��ӌ��
�$M\k�x¦R3�UAP�|�V���Iğ���̟h�	�� sH��2�$hH�����&�cyr*�>���?!����OA@R��8�f�cr�&�aC4��>��i���1��	� Dΰ��v�4=0-W$�?&��@!���hi�˓&��!�Se�O��yO>�+O�	z�Aڙ����C\0pVT;v��O��$�Ot��O�<��X���	�ez`K�D��E��<R3�Ӻ/��I,�Ms�2-�>y��i�h�Dy��iB�&A	;��Q@�F67�t�D�21\7m4?Y�m�}���O3��x��YX�' �H��3$}�D�� ��kf�����+ozPpfȒo1��'%�8	�' i�iQV"��G>Ja�ħ�$R�ܨ  �/Q�$�p!!уE`�=��O�-�H�t� 	.j�`e�٪Iݶx�0��F�~a(�Ԍօͫ{�^���#Լzzd�b�(FqZh�v*j}�fŃ:"�x2���o�f ӲfBA��"nV��m� ���k���:�|��"o�W��$�I�l�Ԝ��J�5�.��J���1�W��&�9��m�C�D"2��B>����AI�vDt���eb���㦍��ӟ���䟐y�O���?9�'�Ҥ��Չ�C;&\�i�}��Q�wi�L�yR�'���'�4]��CA����cI</�<0�7-|�t���O�!�'��	şP'���t�P��%��J1���[|��T��=���!��?���?AO?�&d�)C�Z�)���\ӈ���x�A�'��	���&�H�I���{�ٌ	����`@CLX��!F
�Aw��	E���	�P��ş�'?a �Of����L"c\�d���P�J�a�۴���O,�O�$�O�ɀ�]�9 ޅb��+�5�0�@�.�yr�'��'���p-�O� �KGh@p������D�6I�6��O��O����OV��2`:�I=p��xe�0D���k!$�.s�6��O������d�O0}�O2�'���C�ΰ���+i��$X1o�m�jO�D�O&����6��r�Ġ�&V�Q
a"�j+���T'�ʦ��'+u��	��M����?9���?��_�����V�*��-KЀ]0I�ph'm�2�MC��?�'�S�?QN>.�jL���i��5�'�@�b>�4OO�x64�1ڴ�?�c�i��'m��'������<��U����
����5aF��8�l�le�?1.�]b�>OX��^I�^	rd�Y�T���i���B�Z�n���,��ӟp�I���Ĺ<���~�G��@��T5Ė�(X�=aTM�&��'�� S��'��`�'���'�2/��q��p��,�6��0�9j�F7�O��F}^����J�i��iV�I<t,�� '��\��!ZrI�>A���<	���<���?������8-'n,��G �2�~��g����6�M}�]�D�	s��ş@��?Tr��򒊃�g��C
�~�ȩ�b��T���w�P����T��J����:mB�SƏ)�B�AV�X��M{(ON�(���OL��7X� ���-�$ �6o׬	5P�@��א_��#�'�2�'M�.��j���'�$�C��B�Mµ�M���UwӪ�$,���O��D�Qؐ����I����\����6V���3&�t����OLM)15O��Nz�$�'�"�'���fBY̺)@���:?�d@��g7��O���ܑ\�F����n�qC�$ϲe��1D%ߑN�j�nZ�Wl���� ڴ�?���?��`G��qw�$0f��_�4�"⋣SY�7ͮ<���?�ß��Q>� �c�N�;E��ՈLk���5�$I��i�B�zӮ���OV���O�T'��'R�5)��O)H�:i���v��o��D�	�x%�擘r������j��F6�A;�Eр}F$`�����M����?��?��xʟ���<B2����%*��!�Bg�5��7-�O��O:����!��$�O|���O�dJ�lU�,�0䂀t`��2o��������H<�O�ɧu7��|f�{"��mt`Xc$�ܒ�ē�?0�AF~r�'I��OJ�-� �Яږ*��`(w&]�S|��U�<������?y���~R���+4B�ʐ	�b�j��ߖ�Mˀj��*�̜�'m���dS�h�'7o0�K��+;�E�Ao�s �Ao�����b��?Y,O$���im0\���t�|öO+�8Ł!�<?	��?q�������O�U{��S�J�U���3�1p��y�?�����ϥLv�'�R�0��v!��9[-��	�F��M���?��D���|��?����df�H�.�X��'L�r	;v�Nt����'tV�����!��\|��"QO�����i"]+�[���I���	�|��kyZw�f��g�_�P����"D/���4�?�)O��2��i>]�Äi�rd�Ee��Tj�:F��lS�i�ǰi�rAc���O����O�e$��'!��Ч��{��ٱ6�ngL�n����I��X%��S�D)8�5����K��2�`��F�؃!=���i���'�2�'��)J���C%Y3-�dYB )ՕUp"c�j��O��i���$�O���O�$6k 6	.t�)�ɪ~�:��.¦	�����BM<�O�ɧu��^/d�HM�����H��|IMX2���?Yd�E�<���?�����3� �|JW�U(!ja+���|�@MQ&�i,O��D�O�O��Ӻ�@8Y����U��'у�̦���"	KT��?���*,O"��<}!��³��.+�}X1�ɵ1�V6m�O��3���t�'�1(شdA�D��n��Rx�	�� p���;O���O����Q�5����O�Dc�E��UG��g���a O֦	�	u�	^y�O,r�~J�� p���@��E*3�Q�w'�Φ=�	�L��	�@�ɻ��I�O���Ok,J�?d�t šK�2/��P�Y�`.�'d��L��b�s�֝�{6$�ӂԋbp�h�c��
H�69{��$�Or�oҟ��	˟��I�����fTKTfJ� ��w"0$֔�ɓ�i��'�pу�O���ɐ%f*�nؐ8�>I)˂H#DQc�j�t뛆�'�f7��O���OP��l}�T�$	-YP��A�s���Ua)e���M��T�<����Ĭ|j@œ�|*��'�*�b��X%O:�"��t6e1ӵi "�'�b�'�������O�Ɏo�)�b��-�����ի}B7�<���]��Γr|i͓�?i���?�֨�#M�h�Ӎ(�tZDW�/����'�J�>�*O��d�<������0�J@5B8bg�9���GĦ���K��	�X&��Iş����h�s��X���C�*[В��1�F(�
6-MY}�]�T��^y��'rB�'HZ�3��]e%��hIC���yB� 
.T2�'z�'��DU>��Om:��3F�bT,�1��vE�yܴ��d�O��?A��?�� �a}2��8Z����(�.�T�4��	��d�	����N|��Q?���8Z�V���p>Y� /!.�T��z����<���?�f3��̓�?���B��)�3� :A��XQf�L4�Z�PT�iYR�'4Rhҟ'�R	�~����?���6�Y��A��4e���G��q�@\B[��������I�����d�?W�;Z��� D�4��y�6J�M"���<a��Iޛ6�'J��'����>��sy�\�3o�5պ��AI�M�`�n�ޟ����wJ牍��9O�˧gB0��Lq�\�D��	F�|}�e`�3c2��lП�*ٴ�?Y���?��-&��@y�Z��\�r�ٟ&�<p�!S�,�b6���[��O�����H�����O.�Rl��c�Y;D�z�+��PtH6��O|���O��d�I}b[�d�	~?Q�ӅU���
�KW&l<�b/��m�I[yB�� �y"��4�'�r�'�.��sM�,D8�mQ��j�4�H�jsӬ��O���'��IΟ8�'�Zc!�Rc��0S*\��ƭW�� �O|�2O�@��)�O
���O��d����U��Ǔ�W�$�s׭@Q ��#1�i������O6��?��?Q�OS���S�+dB���U�W���̓v�������?����?��'����|z����fF
���(���ѦY�'32V�\�Iӟ�������a�����"κ|��v��3���`�O��d�O�� κ[.� �OZc�@0X`�<HpP�@�@<����ٴ�?�)O����O��ā	�i>7�S�`�
�r�'��8����~��V�'c�����yB�'),�'�?���?�V��[�ȡNS�3� d��
Z�_��	Ο�����,��b����y�۟\yP!�P�h�=;�,�~+�ك �i��䑜'}re�|���O����O~�ԧu������dD0.�����N��M���?���@�'��S�4P�7mŭ	\x�H� w�΀0f�N"���';7M�O����O��d`}b\���`�^ˬl��.ެO{��pg㎫�M�N�I~�R�0�OL���O��N�� ��G bM�h"['�87��O����O����g}�U�L��K?1�� G����锓E�q��_�a�V��i��Γ�?����?a��"a��	��0�eR�J��!؛6�'�rl�>A*O����<I���5��y#�ɡgW=~�*�F[V}���y��@�%���'^��'����uw�!Y��!��1y�`�h�,�M�T�8�'�X�<��͟@�	�w桫T���wb�,#PG	��Mc��y�l��i���	����I�?)�O;�擛����M\�*���&�d6��<I����O���OI�bT��(ѦʏV�,�!�X�eNeiE�4mlb�'�r�'���[����~
���2��!tp�QU�[�,ٴ��1j�Φ���jy��'�R�':t��O��Ic�(���	O( �dx�Ɔ��6m�O��M�P-��O.\�Of��'��B>GPl!r�+�$,1F�s�Cܷ=����?����?�Zc��7���?p6D�e��ɫ�m\�P´�"'�{Ӛ|3@3O���O��)�Iџ ���ҮO�ь�أ"EԖ9�R�׆��
����'U���yr�|W>�Cp�y��P�c�ĥD_���`χ]�}q��iIZ�6�'=��')2�>�)O�؁�"��@;!�X5O�DPy��Z�y��|���Hy�W>�Pfh>��	`��J�N�
R�e�G���^��۴�?��?1�J{��Jyr�'���$���$�\�d�`⭘�7���'��I�`��牭	��ȟ���П q�%;`�I��%��v��U�� ܛ�Mk��?1�^���'�RY���i�]��B�:МuZ�j�: ���Ƽ>��A�<���?����?	����Ӻ�A�[9 ���pO5M�����L���0�O�˓�?�)O��$�O�DJ>>�4�X�IυOhD�Z N�q0$��=O�si�OV��Ob˧��I�|J���b�F�R#��'3e�䛐�����'�bW���蟴�	����	#;�|@o�*��|�D�-vV��`'^ǟt�I�p�	4�u�'�rC�~���� >i���!��-Cg=9{ft���i��Q���I͟��I��	ݟ��ӺFľodB�Iv+�.gg$M�c�i�R�'7�� �'w��~����?���iTJ�y�$�I�8ђ#҈W3���x��'�RlH��y��|�ӟ���%�Ż^�ܤ�6C޼4�85�a�iA�I��'�R�y����Or�$�O�<�'@����;�p�h�XX.P��4�?���c]h@�������i!}_��D�*_��0�W�2N��y �,�Ms��j��f�'bb�'��b?�d�O^��7��07¼-ȱ$�	ݦaz�H�)J0�x��$�\�O����'��L�$�݁�H��t=�<"�N%/�6��O���OD���]��?1�'��T)bo�z�@�Q��z�4��=NN��U�Γ�?1���?�R䉷,�(1�U=~�6Q@S1K����'FB 9��ON��"��Ƅ����T�D�;!L
�Sbm�f[�0����ɟPc�d���Iן���J�I�q���Dތ+'ņ�#����!��ɟ($����ɟ�B+�-8����Wd��K��Ta���C�\��	��	ԟ������&?*�O���0c�k�4AD*��n�Zt)�O$���OޒO&���O
���T�$[D�I�8����\wɞ騂 ��y��'!��'�� ��O��	�2iЙ	H�.s��IEn�9s�6�O �O��$�O��n�O��'��5sD���F�DT)�dR�a$�H"ߴ�?a��U�d���?)�X?��	˟��I7G��q�U�ݱPV���@\2��N<Q��?I�-�?N>)�O�Z�3DJޔIhx��ME�!���4y�4��?��i�r�'W��'z�E���KaU�L����W�ˋ9�:�n����	4'�x��f�	^�$f��M�@�8�]�F�ؘ��,��]���M���?����?�t��b��� �E�)������ZLh��ܴ��������)�_���O� XTOC�t,�Y�	�J��XA䦕��şD�Iڟ ��}��'���]�H>�3�%G�]��D	��GZ���|�Ý;��F�y��'���5֩�C)��c���R�������MS���?Yu�D�Ot�Ok�A7W���;��͝�D�����	�;h��>w(���p�	˟���Ÿ�%8��[୅�Y�t�H�i��Od�-ړ�~ro���b����j1P�Q��M��6s�MΓ�?����?�L~ʁ=�b�hDoP-{.|Q�I�$ �,�@W�$��B�'
�I֟ȢGM'AP$�	���C1j,�Rd�1H+���ɟ<����x[w����(�Iϟx�d�%f�@�+�d�,]ʼ�E�ϱ�M�����?�/O~���x�-��sO���v�J/C��%rE�Q��M���?� �<�C���П(��ȟ�9��҇g8����%/�<�U�ݤ�M�(O*˓8��(������Y��UX��Q5���:���6�M�ÄG�?����?!���?���?����?��$�W�zZ6ǖ�z
)�c懽@\���'��	�L�"<�'?�dn54F 9eP� �<���?v�6��Onǟ��IݟP�ɝ�ē�?�3B�'nt�yt"[�(y��`$��p��6�C�O��+C���I��q�_�S������>������M����?q��?q��$�Oz�	�#�n� O�	�Ҹ����(ʒc���P�n�x@2}�p��՟��	�[�@$p�i�89F��k�(��	�D��4�?�N�'"�' ɧ5��M�!>�iI����5�H3`�'=&t��'r
�
�'MR�'g~�����<w���I�65��4h�L��UɊ}B�'F�'eR�'�b�`��4OfU"Y8P`����bY��y����y�'��'N�O��蠑{�d4�����$�<)ѶO���+�D�O���I#=L�I�
��2�U�]�fIc ��0�|�P�'Cr�'$�!8��l���'����DX���Ĥ�4� �BT�h�@�d)���OB��X���'���Х�U]w$Y"#�Ż5�X��4�?	�4��H��?�[?��������	]%jxYb�'>�� 4��#Z�E�N<����?�gLL�'��)݇}"	o�+%h>
d��"!�N���y��'��6-�O��D�O��$IP~2�ٽGn��G*	V\+�m��M����?���@���i�?&1�V�!w`9��"D�u�<
�+�M;���?���?a���?�.O�'c,ꕊ���Lp�m���W�B�:V^��yd�<��|zE ��<��-��D�ᧇ�0�$��hZ��|���i�'B�'�O6�'�?���>[4x �(,�x�ґ�ɇXg�OJ���6O��+>O����O2��q����!����\�sea%Mmߟ0��Uy�h�~j����?��� qh�{P5c����1�x2��iǤ��'#R�'��O#��%�֨�d�F�I�
!����>H���'���'���'H�'���OnxKu.#�x�:�X,]8��*�iVP8�kȰ�yr�'��'G�O-���]GLܚ��eM�`�S8f�ꓡ?a�����?i�{B�׬����M���T��0bՒ\;��	��I��2J|RbS?��ɭ޶HC����C�^�r͂X=�޴�?�M>1��?����|�OH����j/YVYHÁ��:Mo�������t���	蟀p�����O��[�Yd@)#F(6�pƈ�".�4'�h�I���,u/�<��4?��R�N��j̘��E�tmBo�//5*��	ݟ���؟����P��Yy��+� �|���+H�<��0C\�k��qQ�i�Y����c3��|����}6�,Q|`%p&�$3*�[ABv�����E��̟��	��ԀM<)�Oo��cfMA�>�L��sH�?^��4O=�������yl��yr�'��
a�Bs��)�oK&<z�\��,v�
�$�O��D�O�˓��i�O��I,\V�!������\j���S��89��d��K��F�<����?9��+�|�@���sfnX���ҕn�B�
�i�r�'��b���In�i�E:)ˆ1�&�sg�9n`�ã��>����<)����<����?������n}��Sp���{�DYqs@צL�7�s쓹?�L>1��?Q�k��-��%�e�/�|�;F� B햀�%	&�Γ�?���?�M~b�>���r�5/|�����$�rt��\�p��ϟd%�t��ϟl�M�>y�>Q�)Ї����,�f�Ixs�$�O ��O`�&>�訟b�$�wאe����\׾A���8!^xinZ��&���	��!��1��
O/����Ȏ��uC��8w�7�O��� ���O�)�O��'��#�79!6�Β�� �aX�����?����?9#��<1O>��O��|���^�W� ���*s4]:ܴp��,��?)u�i���'0�']��Ӻ�(����7(�&���h�DKߦ���ן02u�t%��O�y�۴}�°���vj���C�`ꪴm�֟x��4�?���?����	\y���T雔��K5�u)�_<1�h6MS�!��IPyrU>)� J{>U��D'Z�am��+�BÆ�[@��-�ش�?i���?)��y��iyB�'����96�~)��I�h�H��GӘv��ny�	�y2������'Tr�'m�ї��y{n�I�<:,����Ӱ�d�O���'��ޟ�'�Zc����t�,Yڤ��n!4u>9�O2��7O�\R6O���O��d0��+�7�l�#��ӧW&Dx(4�
9�M��V�\�'�RZ�X��ǟ�	�B�b���ʇ�6(H�%E�" 6���aq��p�l�������E U���18 �^�
�qJ��G�I0���I@6.���b��DTy�b��k���A�e�&[n�R�J�}XnH�NO.N�a�rd�_�@��W�&=���G�8�)�䉖�t�2Î����H���V<u�E�dFD��j�Q���nB���,\?\�Dmࠊ:��`Z��Mtc�����#(�3+4�p��N(h���Pc���
��s�
yx��"&�܇]\�"�,ȪU�"%;QO.��z�@�),ڪ����}�N=Y��P3lv�p3c
E�{���BRh��$Z���'?4a��&�$)
�(��~"� ��'�"OX�:�,���d׉DN�ԧ�i�|"A�!P ���ę8��A�N�V�DC(KW�͂Ǩ�Et�E�䇜�QI�-��)�}�8 36媞����/�O���)�'�?1u坢T{Jx+���<�a�e#Tf�<�#��@��T�T�L4-{����a����D�#1 �CG 8�̓u�H���'a"�'� ��O�'�P����,���
�,Ԣ�B&֦(�ӎ�+��	"����5�$�3���k����I-,��n�"s�ձwG*��dK.M�V����L>�3$�+��4 �C��bev���Շ�?)�O��P����	�x]��ԏ������+ZGnB�I!`�f�E$�?*��DÂBэ!Ed� ����'���+w�X2����
���&�<*Q�}JFËŦQ����L�	|yR�'�23�����Z=l6q[�Ɂ�>NRH2�k;p�vmb1��Q��x� �)<O���򅁃T\���3���N� }�T&�976ƀI4#����G�><OȌI�C��t?�v��vʥa�,�6��'&ў��?���U1j�&X�C���ճ�-�O�<ᇤ4  �Y�ꉬT�j�{%w�+>�	yy��+]T|��?!�Lö~����arT�ӷ拞�?i/O��D�O��:��	pG�E���'X�9[�o�STF����3F��E�Ǔ]9��`�l�8g�Y��O��[����ո#oX86� Ԃ��'uf<[���?)O�,{E��8����0h*<|�P��$|O�ݲ��X+Y�(c�ɇ(r�q�OR m��+�$����:
�,�q�@DH��I[����8��֣
T� 9�v�9���R"OEᄫ0y��i�)4��L�6"O�a˱GQ�t$��cʏGOf8b�"Oj���*MH�u�w'�k�FD�"OԼ9��]� ���y���o�U�4"O���e$=zl��Ú)@��XcP"O<$��A5��yiV#]�}z$(��"O�4*Q Z)efb`��"C:1f~$3�"Op�YeJ��}!Ya��>`O��a"OhpJ6�
a����"�м�U[v"Oܩ���	;�(Q��<
�$�[ "O0]�Q�@�9�R�;� �~覤�A"ORqu�[�>6��k��H�T<I&"O� ����Lڔya�)H��űU����"OHh��D�F*�P�FMc�� w"O� Q��7
Ra�5��{	�ٛ�"O�|PK�'Y]�	0I
�
�L|�"O �UlW9Nz��eh����u"Or���t�N c֤�v�p�"O�`BH�-|�Yʥ.B'����"OH���� t�TpP.	����ڱ"O�哰�pd�(cӌ����A�"O,�PdmN����rb��[��� �"O<qô��)��\[dQ�t�4�)�"O؍@��ʖns�4I1%ø^*�8�"O����Ǚ�k����nìdad��"O��3ԭ� @�X-`ToX�pQb-qG"O 8YR��N9:�@W�`I|-jS"O)R"�x&XPq���L9Ll��"O���b�D6�Ƙ�o�81zlB�"O��Ѵ@ѡu���w$V'Fء�"O`eYPE˽5@r��w_iިbg"O�Mj���#_@��7`)O މY"O���5j���z��Ae���^�bp"O~��c���
�
�QD.U��{�"OLh�E#P�t��CΉC��b�"O��Swn��A��Ls��K�7��@"O��R�AG�["(��E$(-�1p"O��{�m�.z���q5O�KƄ�"O��	�I.�1��@ەm��U�"O"�c���IĂ��pB��]�H�2d"O4MX��B���t�şn}v8hc"Oj�DыS0VHQc��IvB���"O�x(�?FRmw��?uiX��"O��D�H1�<aF@>h`�*b*Onqye��:0oz��$�X�$Sp�j�'�b ��IƱK�vIקO��=b�'}"��8-�AЦ���I,����ē:u(D�d��rr:4�u��11B���@	�yBMϭߪ��t�ÙT��Tö�'}����p�KL�S��?q�-�)y�) ӎץ!yX��	�t�<�&.ͺ1�9	k�\t.��fUv?���H�\��|R"/o6�	�aE�R� �(��٢�p>�D�-c��䙻@0&�K�$�7��ے�ҦN�!���(,���C��[�KMҩh����Q�P�!��*����cC'���9`�կ��"O�p˔EH,�5@d�ǫK����H�@���}���'����	��5]��*�M��QC�̲�'���c -7X�0%��NrJ:�'x��b�!�O�ak��#�$���������'cDhB�����"p�ҼQ�>qk���04�N�T,!D��w��(q)@M�"�_�'?h1kU(5ʓR�B�P���5	'��KU���G9o�zB�I�P�B��5���#�\eP����*�O?�DE3uzfL�w�@�d�l�#�'5z:!�$�����#L0M|�s��чh��d_l�'6�$��{��V9`Y��/<	:�#@��p>��38���Ie�X*3[
�� %`X�8Ҝ�O��@�`9LOĈ+�G@�|(�e�e�2C�8����	Zj�5����'0�]�r�F�V&|Xc��^�`@b
�'���#V/H�I��
j�Qƴ�ۉ��Y�$�6#|Z5�
0M������x����I�<qc�Wʾx��Lǜf�H�#�SOyb�
1{�OQ>ɪ���V#<Xj���C?x��B0D�d`� T�.Ð��HQ���7K-���LY����p�SI��A�\���H�*L@O�Y��i�6De��(��73]8��%��$/�!�� ���T(r�(�� ˝H����S"O�M�'��{����1���8f"O`���恋|���7�ڳ7��;�"O��'ø6B����g�"I
�����'J���t�d]�g.���s��+ھ,@��S9�!�$�8�ò"�	�&m�e�E�1�'�6M�����L�
�j��`�9t�|e#
9NC!�$���SR�V z��h�VM]�,D�O����)OK�BH�ʲ��-(\���K^2��x!A�P�X�ף°DJ�1�E��u�JO�e��Lӄ7�"���b�&���2S�'�2��A���^�X�BA��=��Q	��I�w�!�¢3!��#A4�����J�n�!�dK/�$�� S��#����5�!�D@�7<�r1+��4Ih3���2�!�dՒT~P�4ϛr��ԏ�=�!�d�����kPڌxf���D�G�!�dK=R9��x� �=@GJM2�^#V�!�J�nZ���CV�#B���&ͿC!�d�C@}@�0y�\�!tN�p�!���*�=�䎓u���#S�!��^4T�Du�V��C֐`"��^�!���'TA��)Wǟ�B^��!کi�!���%L���`S�n�҄����\�!��N�H@�R�����(�Z,m�!��ά!ҡ@U-5��TГNL>'�!�$AH> ��&g�E[�*h
�'$�9`��I��L���_���	
�'��B��sx`gd�9Y�<���'�z3v���B�hb�.E6Pxͪ
�'��+�LU��.�[6l�M�,(�	�'�J��S��C 8�!6��1`��Q�'�XM˅b��!�L�"6��wB6d��';ưAu��cD��!6`ω
��'����a��"��u�� �\a��'����GeNzhRR�X$)�*|�'�m���,Q�y���LBI"�'c���$,�\��@ck�~�f3�'M�M�#OY;QX�R�K�n�zh�'�H);�U�!�@/��d�����'�x�P,�������L�JQ;D��+�B�ˑ������<ai�.N�H�*�5�X�"A	WyR#�,�<�"	�J������ �]���Y���'I���ʭ*���j���O�	���i��������n�HN�X��$3\OnIr�)I�	�$�'�&eCS�_�gp��(�H^�}c����°M�����8§G� �;��� D`��x@�A<&q���=aU �<y�2���K�O!8!�R�5L�I�QKB��	p��¦q
7��;-9�')�#}J�ʎ�m�ɫ7j�|�`ݙew��蚦@��~��Ɇ��Ӫ��,'�t*я�)A@n�񱍟�B��\�����cc=a��]��	�PL��#�S�nw�Bd��t������U8�.���� �|YB�a�K�\��'}ם�"M���S����������U��,�m��	��y*=�MyÉ\2G:�X`#�_�%)�����O��%v��X�*?
�m;ǁ<}2<�l�P2h��F7x`�
f��0R�'L��d���X�\�#H�2=���3�[1H�f�F�7y
xcW��{��%�(�F�WR��O��8�X�j�������R�p$�W�	��@���@ |�ecu��&����ѕU+�r�eE?^��"Cn�ly����h���	_�f���J	 ��]*BfR"F�6�ό1rR(#����MH ʘ2��O��p"���n��z-r���(͐'8)D�P�Q�R�O��h���<v�2!i'��_�.��P霶X���a�$�6�<q���S�KqO�N��z�ʓ�LK��*�!��0?�^��	��lK4 ��:7�݀q��(�cN�QN�Eqˎ3���'"�2�����m��
K�%ҡ:���Ԣ9��r���
5۬��jY��?��8T��	�'�* ���g-I��vB�ɒ,���玞I��J��F"`ϒ��ߌ1n�Xr�lʍd�h% �$ٲl#?�� J@z�M���l�dڨI�za8�"O� �e��&��ʵNA�����
��6M��9�(j�ϲPPZ�g�'�,h�h̚L�� sꐖ`hؙz�6&�����ByYK�N�}(�i����A��(�O��t��Ն�I�`b�87�Q�	��ڇ�ӛ
-�"?�6�'��ep`3#H	�����:��A�ȓz�,�cQͥv
�I���[,K���ȓ��(A �-�* x�G�0xe��ȓC!�}����<X�y!ܩ��1�ȓ/�~���A6_p��d��K|��
d88ӦA�p�'hތUu�`��B����6*=�`�Pd�]�fx��'��E��iV������<ꀆ�i��йfD�-8�p,zWJ� �L��( ���UIɏVd*bR��AJN̆�@M�� �XB��T�J�e]4��ȓS-���PN�0��IЃ�
\D�X�ȓ;7�EGÑ�M��`��ǽzx���&�t�h���1�P8 / "z��=Up��/�r�Vb@�b~,��0~�f�J7V�����$r�Єȓ���q��7`�H�{��(�����I����r����sm��ȓ7n�`Xa�֟G�.��R�"�>	�ȓ<�V�P��&��8r����h��ՅȓY^$����в��b�Bжw\���ݺx��D
tIr��@X}�q��|
l3!�J✄��BG�)�ȓKk�D	ɑ	n�R�rE�9fb�ȓS�}A�l@4t�V�4�YR�����F&a!�B����Ҽ6o��� ɠ��&�Կ}�t�q�=d.��ȓ1�1��H��P ǃ��(��l��%d)�Ct>!a�B�qJ~C��1(��79!�P,8ЬC�r��ȓLX��9`*��>#�|�af��U`X�ȓp�����b�.��h���_�	���ȓGh���U/76rI�2"O;a��T����ק"l�x�'ؼWՒ��ȓ^T�(�#�`����wH
��ȓb�(C�ȁ#HCt�ӥ�-�E��E��:��N|���'SǴن��؈��)�0�TK'��2sr�h�ȓ�%17�4�;R�\0ea�|������e�+���2���*'�X�ȓ_n��"ѩm,�B��+u�,ه�='ڡ�u�N3?��y����=b��ȓjj$V-�!K���3$lْ'�-�ȓY<�I��A�9=���a�E��ȓ����u��21gF�0�S ;�L��F��DH�B��k����E�����ȓX#Z�1�K 0�� (.D��ȓn�h�l��!O�9��!�,:��	��/Ɛ�ע4\�"�� �Cgڤ���6����"J ��fΘA!���]�@���iD6�l��2�ռ^��y��f�CV䁣]2܊�+K<��P�ȓ~��GI��?|�T��r��i�ȓ9��L�$��	4�9F��	"�Q��Y��rT�S�
� �񤈜0[�\l��� �¤�2�U��a\"�ȓf���I���]���0���y���<@8X`R�J���Cߴ�y���'g�܅���0=�~	kc#�y
� Ȅ�ܸz�d���� &�$��"OP	�%�#!�&)x���	Q}� "�"Oԥ�a@^U$x3��_a�L	�"O�T�ը�^�]K��D�=}@��"O(�� i�+ �*��T�`4��"OrE��R//4�y2ũ�=��@p�"Oި0 �&[p�7)	4Z��B"O\	+��FZ�(!K���+X�Y˲"OD<s��L�\>L����>��5"Om	Ҩ�#i-Ԕ���(W��R"O�)����?xz�ܡ%@�8�b�[�"O��{QmL1t���8��K�kİ$"OFe	��
z:Y�����Ve� "ONk�H�..��&.��
��T��"O�![�鐧,	T�M�8#DA��"O�Y��=L 
�*7��0
��a�"O��1&M�7&լ�9aD
�X3"O>8�兇��9���Ն'd�q�"O��)��� P8i)C�%!�Dh��"O��'*{nhVi߫r����""O PaACX�eޢQ��O��{�"O.0H���G(<x�5��&I^�Y�"O\MX�\>@"�i)g/Qx�c2"Oh ڂ,C!s��y���]�v\y�"O��! ��Y��X���5]��ab"OL*��2u��E �M=,Vc"O�q�G��q�S�懛XĤ�:"OvQjbM�r�\ �Y=��M�"O=�I�&'����sh���TAse"O��`�YW�� �ƈ"m��{q"O�X�7]\ڴ�h���<b��q"O
`9P�ΜLv����Q3p�`�"OJ�*���'{v䀘1�L?|D@XB"Op��BhJ�gSD�-�4&>�9pF"O�|X� չ H�]����1%FУ�"O�K����i"J�r��\�l�"Ov4�p9E��A©��uV4��"O,�g<!�ݛ֎Y:f��"O&�P�(�mA`鹆L��(����"O��з���*�
����#V4��0F"O\m��G�?3���J!Q���'�y�Z6�x�"$�X2 � ���K/�y� G�`���� ��v�iC#�"�y�� L��U/�=y���9T_��yr*JTLZ �ѦK�vMx�!E���y�A#bCҡq6��]�0�j����0=��«��#�u��N�!W$*����)�y�N�l5r�KՖ/v��A�yr/��Z��K1n�7��u��$݆�yB�2`�傡�.
6ػ6��y�f11݄]�uB�mVʠ��` ��y�������7-��l�&@&I��yr�A�y��H�P�1)*�
�&���y����u0�yFh�8rV�0A��C�y��
|7B%1��q
u����=�yBdK�N7,�b�ǋ�c憤p��8�y$Y ����!b{�8�X��y��L��@���_�Rc.T�v%/D�<ADG�eg��+�璁6� {@�'D�䀦@dy(�S�*�>�0!W�$D�j��@�42d� C]����<D� +�á��|���ȧ!���"�g<D��H�%��u�rԂ<���0D������HY>���g�8|�ʤ�G0D�� ��z2���q!��PL�q&"O^(��J�+;�D�[2��,J�M��"O�y�f�k�^���N(X+���5"O����cL�u���F �L��"O���bM�IJ�\�$��(2����"O<���V0	W�X`'�  �X�"O]Ӵo��B|�D�B!!�Xxj�"O�`�#�!}"V��X5�-�R"O� 6�I�S��`@�­TzB`�"O@��6M��N�Ȝ(�"Jt� �"O쉒�AI:�0`ʑk̭
SΉ�3"O�l"���+,�,<���C�oDxtp�"O )���8R&*�hi)R5�"Od-Z�N`�H� 4)ȹ<6�\�G"O\ɣ7�<�<0Q��&���"O�0� �N9k���w��(k�b
"O��rC�9@
�5KB윣l��k�"O���F6)�@rd�	*�A�"Or0
rf� H��<��!	*5���7"O��  �U��<�P�m�:2Ż�"O8�Ԁӑ-�|풡�ћ&�b�AQ"O>���f�!�J�k�&��F���h�"O q��C�"�b�� ��#r��YY�"O^\jm�s|�� �P�$<j5á�'��'�V�ZD*�活%�ڵG�n ��'�l�!��Ӣ@�Hy��#E�2
�'�<9�#���Z��y!�"�2��	�'���V"�Hӷn�.N�P��'�(�o�*����d	�T����'�x�q'J�sy�@�#�� y��'� p�� �j2<��s���P8�	�'�4sC	x�NP�������'��:e��6M��� ��@dr�'(�\+�N�M0�:禚>'�f��	�'�:,!�!D�C� 4$]?�
aI<!��O�v�0(@3����P"���n�<)���D�܃�o!O���(i�<!��`�(�!_*����e�a�<)Q�Z�̲y�
��]Ԉ7n\y�<)�g,Nn<���ҭT<
��/�x�<�v��e�F�*��Af/�|3���<��Ƕ:�l0y6΁�{��C 2OȔ���IB~�h�!*��Dc�"O��a�I�o�� 6AH*3̲i��"O�
��B@�2L�WL19iZX�"O0l�e�&K.�<�@�J��qa�"O ��"�[*YQ>Xh��@�I�Ti�"O��ғ� S�hY�Ĉ���I3�"O����.2����E�t��ũ�"O�*%��Zf�!3坔o��P�&"O�T+n[�hAx1����LȂ8��"Ov��aGĒ8�hq���@ .��`�e"O"P ��O19s����N�.Mv���"O&Ef�ş�f�{�M]x�v5"O
�J�cKB��<2��F*<nd�+�"Obi�u��.�d:3�� �N��"OV�p�D�!�nd��IWH ����'���w� ��dޒ!����͸U�!��ZO�~L3D	/\����<�!򤑂Q��<;%�Y��hXdf�Nb!�P�N��'̀O @��/Y"9V!�$N#u�^�@���ޝY"�ȳ5f!��tN&�rgN�,Ί�0$�Q�f[!�dS�[�ba���p�h���"IZ!�� �3�钊� �``6ƽ�'"O<��@ۼ
k�paE͜r
0��"O�"��' [�5�Fn�b�Ĺ'"OJ�1��/_�`+��ɌM�@\(%"Oes%�-:+\d.K�T�:�7"O���ț�u��P�ȑZi�x"O���]�M��!#
$aR,�"O\!�DEL�(e�r�ԉy,�H�c"O0eYgc��Nb��F�.1��1�"O� ��
�(�ڴp�噠a-��0"O��E	ͫDT�WR2$4Y�"O����`[�SF$�Rj "Ip�"Ou���˧'P<��R$I��
`"O�Ufȇ@f�a�W�q�n"O�I2�BYW���8�$�P�"Oa�)�)mޮ�����=K�R� e"O��v�¹�H)��3E�0�:�"OȰc�NՋ:f�����J���i""O�Y��k�(0)��`�-�ЈP�"O�����I��!��@�����"O�Hh& 7]�x�ʜ?u�!*�"O6�3w��6.�ȓ��:;O<�"O*T����&�pq�rmM��y�"O��$U:' ~���֪�Ԉc�"O*-�e�^��AK�"z�J4��"O��C[S�������퐅"O��E�1Vh%8��Ne�^9�"O�@�/��t��y���7-?>�P%"O�i S�Y�#)z�c�$߷W!�]8B"O���r�H�mCiD:��A(�"O� ���,f�iQA�@����5"O���nW���:��N03�8��"OJ����( @S��/%��a"Oha $���!c��K!S	xU#�"OV!� �Fq4A��jPx�
�"O8���5i����`�[2p��L�"O
�RN�
<��=	�Z�r�.��@"O��UHD�-�P`�G\���B"O�U��o�a��Lr�`ȉ9˔i+4"O���W�)����`���Ñ"O���ChοKl��_�ay�%�"O
I��!0�1&��0w�X;�"O��)b��!"����;8���F"O�������h���� �X&ޡ�g"O>��Ǆ��<��dQ��lr�"OZ�Ři�
�P�ΐr��a{$"O��9��!zb��A�;r:P*�"O��	+�	�8)��@\5Al��H�"O0-z�� �D�Q�o��C0N��"O m��%�1�y�e�R0 (��"O����@�(��YS�AZ!� ��"OZ�91��o�� &�IP�q"O0ؐFO��&���Y�+F�diq"O�9��X\a��k�*A5��IB!"Oj!��.�t� 	�&
�s�^D��"O`�F8��#���"n�D"Oܝ�GA֙E=�8����C�jP �"O^�HvƐ��B�׳:�^P""O���P"�%X���A�z���xT"O6T���3��)���P��&�ȓ&����hǻz`=��K��>�>�����dJW�A�ϠD�-P�.'��ȓ]����6jװWt����H���8��ȓB�*��J�:?EKEc�����S�? �Y��\K�v��Ei��Q$h�"O��"D�!��M�f���+�D�P"O���q��8YB(�&�#=�j "O�a�c��80T^�qVV�su:��"O.�� ��t$Kwc�4VZ���"O��
WvB^��×C<�}bT"O��3� ٴ�Yp�S�u3�Y�"O��Ņ�0jF荙|%�܊B"O���I��n�5*C�%vz�`�"O�)8�(�*���j��]�"Op�`"�(4QĤzuL� �.�YV"O$�(�Z����3���r�d��5"O8q��l�F��=2�F�<��i1"OL�k�&M�p����&�1��m1@"O�����ɊhxDA���Ҹ�Җ"O�9�s��t�Y��Վ�x�kW"O�9 �N)8�y��V>�r��"O������K�$h ��.>޸)��"O$XhG�S�)�(��Řs�6E("Oj�q`g�$\�}�)�4C�a"O(Ȁ���;�p5C�fZ928��"O�] �A��J6�|J�$Ph* H�"O�=�Q��C���R�Y�yԝ+A"O���DG��^tB�I��d�!ұ"O���u��EܨA��G.xvQ��"O���q��0JG(�"��Ϗ*��@"O���3�M&���QX��"O����K�&��$��-S'2�6U3�"O8y��*X�`�ҍ_�RTp�"Od�fk2��@9Q.D�x�\@E"O~�:0
F�t�!A1�P�O�J�K�"OD��JϘJ�����6��MU"O�8[DA\�{���*�+�;-���r�"O���ň��w	�m�TK7u0���"OB�X��פHi�����]����"OƁY��ǿe���e�,W�H�"O��T/��&plx�%� �P� 6"O��������8Ѯ�w�nh�"O�"┆'L�*$D�$-��p"O�����=&��r��XP��("�"O���#tF9)%߂>>�ݚ�"O����H�4%���u)܍3$m��"O�,�S!�0N�A
���4�J���"O�".��S& (��^'xԆP��"OBXG��
=��#U�b���P�"O���wjQ=�L��B��l�~�Q"O&%&o��)�n����]�|���"O���gAR��iM;����"Or`��G-P�����b�T�n1yC"O����\,#�9��A8l���
3"O�쒠���M��+��-��m�a"Oژ�)=nhp����T�PH��"O�����7`���(f$an]	�"OLiaM;�P�(t�Z�w�4���"O�]sv�]�u���c��т��]:D"O|�u%J2l�T���W���j�"O���!	��_�T�pL��0x�"On�Y$� fp���9�lj4"OK�4�����,W�$�� ��y�(�73b������Q$F�jw�"�yro_��l����Y2F5�yc��:�yb.IS�|�z'hM�6�؍���V:�y2��&QE�I��^�.z�d�w\�y�3�82',�'1���w��y
� ��ǆ1b	� D��7�H��%"OP��<@��Db�i�J��Se"O2�bF��/)Ԫ����\bm"O�M9�lI,��a�"�	�JH:a"O��3j�-���cB�T��	�"O��:`�5k&y���9 m�"`"O���g��lpyKDkJ4
h�8"O���7
_9-�l-�5�7[Ӹ��r"O�X� �.=ԫ0eW"� ���"OZy��_���&��5�Ԁ��"O,��ϑ0Ő�7�2�A""O�Q�������٠�L��e!"O����MI7Z&���#ꃪ �(|��"O��25D/iS@éQ� ����V"O�)i��E7^�(-���h��;e"O��peb�թŉ�'`c��C"Ot� "�5}��`���}E��g"O!녉�P@R�ڤ��62��c"O���$�C�
:|X�'�sѤ	I&"O�e���]$8E���'�/��Y�w"O.�XS���5`�#�	;B<0[T"Op|�rG�^ך��o�W�Xw"O^ � H�5�*M�P'��p����"OZ�!+�m����ǵ��,�B"OF�!G�����wfτٖYr"OD��%g�F2���#E7z�P"O�Y��]�����5���˺�Y"Oz��%W6S(0x���:�L�X�"OD�[��܄0�"Ġ"�E�n�|`ht"O,葦k�.�Ʃ��`4-μ�h5"O��zQD�/N�j�� �S�^œ�"O����,/r�����f��F"O\�@�$%9��:�M�=�l0�"O�Y�C��,m�x�s��+:�>d`"O�Ī@ G"dB��Wⓣ'��A��"O:���'�usF��s"OFT���� G��!4E�uq�Y�a"O�q*e�<L�V��s����A{�"O�\K�K�1/ZR��Z�i�R�y4"O���N͑@.L��$����MH7"O��Y4↭,8B�aOR �b�{"Oje�R1���)�1Xrt	�"O¨��Sd"��{S�ɕpj��e"O�|�!.�̘��L�	,��F"O������I�"�UK�ibp"O����.F9G�5{#���-�ʐH""OL���b��e������5���B�"O�Iː
�	bdڷ�L��I �"O�� ���z\�BA�C����"O�!qO�H� 8X�j� ;��1"O�t�w��2q���cp�F�y���"O\}�gͅrl��(���;~�p��"O�p��-��#~���E��e���g"O6!� ��+@ t��%�)(u����"O =��/D1]��d$�*k�p��"Ovpu�VW�*���#PY��z�"O\�趢F�V�	�ĵL% ��"ORE�s)��:ϸ�#%�2K��z�"O����W�N,)�d�C��(sp"O�Y��_.Z@���;�l��"O�QY�AZ�^�����P�Tǂ5�2"Odx��a��2��L�6Űh�s"Od�j Ϲ��Yoމf�8�U"Oz���D�.i;R�	�h���	�"O� x�J��3e5�p
4�T�FjVus�"O���$"�
�p8�k�`\��0�"Of���J�޽(�䞛i@2g"O� ��A�7����iA�VZH�"O�͙ �K!��$�:6Gp��"O(�id�ؕkp�mH��k�B���"OT�I�W���H�#DN�l���"O���8N}\�2Fc���� P"OT�8�h�1n����@�À,"O:�pp��;�H��G�A;ь���"O&E*!���L�{� �p�8H�O\�
�,V�:�d="�lݜ  ��� �8D�T�22�28��qin�֭5D�P1�� q>��``�؅waFu�4D��k��S�Zk�H�+�h�"yꧏ3D���c�˛!n�;t�P�9O�\��C7D���OH�N��䙨k���06D�d� A(�BH��b�.,�袦�5�O$�	�Б�g�f���S��5B�6�=���D�OZ���W��XL���6�`�,D�����?� � ��	r�&T�6D�sR��:E,�ٳ'H�y�x���5D�ȩ�aL"Ἐ@Q�]Ȅ>D��BqD������D�e���qv(;D����J_:k��	�T�УB�����#D����4�LP�U�ͬT^˥f�O�C�	�$V��8��{��C'��"��C��,�N��'g�%W��H�ȟcf�B�I{H��g(ǎ>
!��+�-9]lB�Ƀh���z`뛍���Ha.j�`B��4j�u�̋f�iP�	&���[�p·K�CҶ1 3��Ԇ��
% Q��S�"�
K�p�y�'�a~Roɴ*{�M:c��0�$m�>�y��ė$�|!jR��T�D�&�
-�y���8�ҭ���9t0( 6lͦ�y"��6
#�<�V�L�Z�D˶%�3�yr'�gi�t�W��/O��Qd�?��'nz�2��B=$
�괤�F���'Mx��Õ�0��9٤��

,�4��'��]�0�O�;� P��G��}�V� 	�'Wnh�"�5A:��w��t@����'�.	�d��� WG;h'���'����!���A��IC����'�z@��퓄'"ݘA�+龠�.O��d-�Sܧ\	иZ��_isxL�ө͸�r�E�R��ɱ(�"sQD+51��B�I]S8�r�j��` ���l޼
s�C�	�:^��'/�'*�pڐ
H��C�	�D0=(�AD(0i� y�ȯ �zC�IC�T|�"(�6�h����bC�	������QȤ�p��*�*˓�?���S�k��;#����1y�/ϨY��?��I��R]@=;C֕?�(�&G߄HR!�D�(HX��j�/�%����/@!�$��~F��#�����i�*�	}�!�Q3o�eX �O8e&�
����Dp!�ḏ5h�����0!�*�'�Z!�+pm�ٙ�ᜠm��Z��գ;;�"4O�`��D	�� Z�_�[��8�"O~@��h[�=+��R�J�|��EX�"O�93q�(��5�4��x�Du#�"O�"胗V\m�k�Fђ"Oرd��>}���Sge�j�v��"O� R@��E�N����1��x�<!I�"O�I��C	�6�L��&�W�@!�@"O���D�;m��x0%��XѾX�Z���'�2]��G���՝J��C�����=JVO��'�ў�O��𱕊?T��Q��YX~}��'��L�a,��֡{�C!FF^��	�'c�|h�~TA���DH��'a>-RQぱ:��� �/A# ��
�'zy�U�*�"� 1N:���	�'\��V�х/�!"�d�>I�p� ��d�<щ��g��<��K�&���"G��C�'�ў�>�Ri�8d��7d��0�!2D���ԧZ�{zzlb���-�b��$D���d�X.0�\m��I�e�L	�!D�(i0��:=i{R.�Uw`@)�a D��� ��K����E*	<�b7�?ړ�0|��@T�YV<��CII��I�!�vx�p�'@*5Yu�Q�@R^}p�o�#䆼x�'m���A]"�b��S�ȵ!YH��'�xZE�M=�$=�W���b��]�ʓ3~�œv1�����)A�y�ȓ��aN�`���Cə�{�\��KA�� �L�"3�y�b��|8��I�<)��ބ&�N$˱���U[>�y�ቚ6�Q��1F,�rT@\8X�TB��3�΀)EE�W!��Sg��,H3NB�ɝw��5�W
�?��Ͳ@�(FNtB䉽�N�(.�P��՚�.N� V�C�I	�|�a��G�p��C)�'6HC�		)�#�gL��X�bm
yn���o���h���S)S������66�I���l˓�0?�Ҥ���Ƞ��o��B�����Y�'�?�����A�Q�"�I$: �-"�*��'�O�̡K�.W7��#W �>w 8��"O�Lq�o��r �z�O�,!�0�Y�"O�Q8%o��e3f�ۢ(٠;*"�'"O�x�	5 ����c�0?�����'��O�⟤�	�<Q!�ͽt�b�ڧ�)�����F�<QFD}�9hA��XW^Q[��Ix� �'��	�Y8��#Fڇ-r�\�'���^ B�
[$�!yEE�p�*qZ&�����B�	�y���s4�D�r*1��ꁽ�lB�'"�����(g�����ýWY�C�	>�t��A��|�`N��:��C�	�7��K�Ʊ���#U+�pUB�	�4��zHJ�B�h�$ "(C�ɟ�,�x��7ZC4�VJ�t<B�I??5R�x$�"�rW	�gz�B�	�gT���g�^����ˠ5<zB䉬@����"U����Պ	|�B�a1d��{�����dN�nƂB�	_f����C\��d�k�-�Ά��Q4 ��@+ЂI���%�ֲv��H�ȓ]��poM5U����B�91�H���}�u��jZEL���,E9-b̈́ȓ#�EM�_0,��Y�Q�E��x��pHƿM��#�Țq��$��et6���a[j��5+���nI�ȓ��4!�+�9tT�0;�暐Whi��O�,��/�
�N�G�P�kJ�-�ȓ+'�A*).V���t"�k��ȓz�-:g�D�:#Jx#'=FZa�ȓv�&��SB�=D\,X�c�ra��ȓtV� B'��n�t��%�0wҩ��S�? ��
��+6��:#�9��p��|��'U�-�mO3[�(3'�F�AB|P9+On�=�������xq,Һ�$X�P�F|+ў���I�.P�B�o�!]*��� D�$�PC�IPe�8:7�Ρ5�|�*�M�)�C�v�HՉ�e�-4�
�a�
x�C��&�P� �
��-�$�^�^��B�	�MҘB�
a���@TF4h ���0?I���v"(@h%��>X�P�e�T�<�C�1Py��1f9k�9;1�ΟE{ʟdc�(�1C�2%lR[¯�#��%A�F&D���Rϛ<Y3x��4���̤kUO%D��ҡZ?T�AB&GP�e��X��.D���2�Ծ0�H-�QΎ:=DN���%ړ�0<A���+�Z9@P�Œ7!�q�W�[qy�'m�`�ʍ{瘑x� ������'�XX(3e��\�p1�I3hd�����'��Ov���<�A쇫o��P�"�V� �(�sB�m�<	�f��6%D���b�] ��6*�m�<y������BL��
��BJ k�<i@��P�$b�B�^��8*�`�}�'�axCӠm��!���E=�@ek��y"oD��(5ra�ԙ>��qy$�D��hO���,�'
�����P';z�mY7G��+.�G{��'g�A4&ɛfJ� �3IZ�>Y���'�m�b�ǡn�h�#.2|���
�'�Ƭ��Oƽb�l���eЭ*�vh�'	�Ւ��kk�X2�(�.�{	�'�(�J��$|��|re�ڤwĠ�	�'Ʀ��l�Jud ��� i����>�'��	�µ�Ҋš���hU��ß�F{�����@�D��UK�����Ƥ���=D���1�H�*c�pѡ�1nh9e� D�Ի6o�_}�`8s�_�5\���H>D�4Tn^���Xk敒��:4��b�$�&�<�든�+(@��"Eu�<�bJ� 6H����ݤ3S�AXa)z�<���F|x���ȩfHnXJ�&VZ����<	���(]��"å=I�Ր��r�<)򁈼R��s�	SV.u���q�<�l�C#F@�)��fj��s�Q�<�D�4E���PU˂:J�$M�DO�<)��ʚu�E�v��Lp��6��H�<q!��1݌�q�n�*mUTQ�.�G�<�s��U�5�VdY$yﬀ�s��A�<qq�ð&Zdc��+�B���h�<qWk�l*���p�t���;/�Y�<6#��a'`�c�!ЄHB�4@��<)��܌w6�uRE
[=*BI��/y�<1Ɖ��"���A��p���	Dr�<YU��W�4�����˖$�s�<��lׯz���,�$<�t#m�<!E�N(S6 �mN `=�%�j�<���J�s���w�]a�^L9� �@�<	T͔"L_�D9V@F�`���ZG�<A!�O�)���2��A@%FuxO�E�<�7���SPFPgb�]\M��lT~�<�bGJՔ���9t���D�Rx�<Q7�Tl~D�����o�\M��/Rr�<��'I����h�Zh8���X�<u'O�}P3��@�n*Xq��U�<��=.�șz�T^�qqKx�<񃣒:FY�Q�4��.?���D>�D���b"C�R�,E ����d��S�? ����w$� ���nǺq��"O|�[RK���a#��N%|�j!9"O�8�4��wF52��.�-�"O�E*c�L�w�t��4o9F��"OT���O�H�\�s�n�i�RY`�"O�-)�̺I�
@aB��J-�U"O
���mT_�
���aڮD0�"O�驢���d�0�?Iɂ���"Opd s���?�&�����(u�'��	���(��U*!��E�T�N�F$�C��;Jd�Kd�E� v�ܙ��1Z<C䉭m�B�c��4'_� �����B�;[��!d�*i� ��"l݁d���0?���B3@��1�S(�?X꼱��_�<����6��i�d�ML�i!!c�W�<q�)���y��Ι:�~�kpJ��d̓2��(W%s���R�)�8ZR)��^(���K0��q"��Q-�T���=�Uk�]�6�
����g�u�ȓ"򀈷�) ��'��#P���%�؅�[�z(�f� K��ȣ���^j�C��9<���`%E9��@Ru��e��C䉅O��X��'^�Ĩ�7���r������/6�@ӕAF�7,|��w�Ɯ@w�C�G�V�p�⊽VGJ�s-F!L�B�I�f�r Q�T-�<5pS�+�\B�I�[-�1��߬+M$];�K�P2���O���D�. �r5�s!Y�T_�ܪ�?!��^I���h�I�2ET��I,��nq!��V���&Ý
~ ���L�cV�'R�O�"<)c��6f�`!���q��a��T�<A6��-Vh��@͉d*���b�g�<���p�N�ʐ \	;-�@4"Bd�<ɣ�<���.�j��Hu�<��m�=k/�	�a��0�J|���N\�<�o��!�LaB2�$�
���N�<�uL��&'�|�5�Q�rr��jC"�R��P�<i�K_T��ͳ��X�O��J���f�<���M*�D�E�"�8)���`�<�.Ҏ�McA�D8<��Ģ�A�'a��O�FK�1*���4ྕ6l�y��-x��'N:2�������yR��/VѶb�.U�;�\i"_�y�H^9	"�8�d͓1:��Л�y�B�7V�hu�䃏"8p�x7 ��y�$�5H���#m^����aMM��y¡�[;�E��Y�,"us �˓�hO��D5�{w�](����aHx���C�_4�]'�F{��DF΄z���6Y�
�����y"�W@���� �<�\!��?٘'p�H�M��P��
ߔ������hO?%�`	>2 �G�Q�%r� �8�$8�S�O�Hp��ĸ$�40�F��nx��"O�i7JŖELT�ek
�ba��r"O��Pw�K&!�i"�؋pF Y��"O��8�F,ZAc	Y(VA��"O$�y򎂓`ȀC�Ι	�L� �'��D%�, ����mx�rU��0z!�D�	<Ґ��V�
��"KHR�)��6)P��NA�>�0vkM��Q�'[:�S1!D�c�4��Ej!��Y�ߓɘ'XrMp���r\��Ĉ-�
0���?9���I@��*��v�S�t�>@�� --�C�}_ސk�#�5'�r���ـ[��C�)� ���AG$Xz�m��@^���24"O�ċ#隤*���k/]�_���;��:LO�����"<Yh���N�8��F"O�ViX'[�,hb��Gs" �P'�'�I
&h�仢�B�\��*���)O�B�IR`��q�@7!�>�⃺3��B�I#}݈��Q��Bi+p�F�+�B��+2��`��_12<z���PT���I^�'f?y���)�c�9&�*0j�)��0<�2'��a�X��UK��5t^)���VI�<�$o�n�xQ��N�?5�����Jx�t�'b$�	��M�<xhQ'*R�~���	�'m�$X4�A�U��8J�/��tn�T��'�l�GH�'hĐBBME�0�R�'��h�'E d4΅:Whӿ=�b��'���VD�!<l�����[���*�'bF���:�S��F�}�
�'-���U��s�`X R�S=-���Y�����*>�^�����5���:4e��!�d_2~�(�g�3x���y&*I+*�!��+Q�kK��G�F���d"Oh�pዄsl~�qufQ!�� �'���9Ll�y��L�iS����˲:LJC�I�ru��HW�Ϣ ���6��5�C�<p_��b6bߜd1��@�3���d�O�{�&�ZrkE-i��3��}Z���Da��*4l��7����J#>����7����
��e�*Q��6�XI��Ga(��RhX�	��Q(q�`�ȓh���9%n]+s�pu�cO�&4|��ȓ�~lA�AY�@e|�q��u���z�Լ	�� ~�7���t�ȓ4�䁈e�	���w��}N��ȓ\ddkBĔ�8����,DA�a��q,���.�T�! ���v��ȓB�|�ZG	:X8�(V�J hB��%��E{����
�N�8F)׈r����ڛ�y�N!����R��RJ�AX%&�!�y��ʅ �x���1=-�%C0����y�'��jmA�Aͮ2� y��c��y���-��	�gi�.*}��8�!�$ȝ4����#-Q,�Cَ�!� =NȆq!7�ЅV.��!!�P�!�d�
q;�;�7F�Ys�O4�!�#�2KL�w�Z{���ʠ"O�Pg�åe�d�"H��	0�����';�Y"?�`���V�@���!L��^y!�бp'b��"W!1N�j�+R8=�!����iEGIfpR0QQk$z�!���3c܀� ����mq5��	�!��|>6-�s'B�\t !$Jp�!�Q�k(�=�P��'{�9�D�$1�!�dJ�p��( `�B֚i��B�]y��d w{`*r�ʿ+�ށxv���~�ޒO����D-mܤ�׬��JSV;��E'NS!�+n�pƪA�S�0�:�cS%Yo!�H
m����SF�����ԠR[l!�Ӕg��*��ٸC�nM�Ϲo[!�dÙ>���H�j�ۓ�$;�E9�'Dhh�fN+B���R��=0xމ��'z�%k4�P�*�ȱ�E���$�F���'�x˴#�.}~��Cd����H�'�\ex���`>j9S��5d�0�'� �,��vA��j���^h���� <�Z��W�m�J�ې��QF\�W"O���A��QS������`�"O*|)%�/^8��_2�!�"O]�Ԭ�37���hp,�&|�I"O��@��6S��,�MB*&q���"O��� ���X����M�_Il)�"O�e�B�ʮB�q��#�98����'�'ў��J�'O�����-;�9�r�
�s���X	�'ZDѨ�oӳ0�N�j.A)��[	�'�~|P')�k��< ���6&����']<�U҆K��D��/��آ�'SJ�����g�`x��������'�I�F)1^�x-��J���*�'d-
��W�-�(2��IL����'�(���+M,^ S7��/q��	�'%(z��%/����v��8n9��'��}(�GĖ{�y��kщ����'yp�c�N1��	J�� *q�Z@i�'Y�\(Ӌׇb�p�b"C�}��� �'�;a�Q$yf��@��?r3���'۬��P`�;xe��	t�,g. Ě�'������Yb�y�é���z�B�'?ax�Aҭ\ x���6�~��K�"�y"��V����s)�dPvkB��yR�Nyr��w�[CZ�P6�� ��O��D�Ob>E`@����c��I;Iڼ\��-D���f�[��p �BՕʀdaB++D��)"�-2 :5���f�5��'D�h@e�ΔZ�>U"�ǥZ���!��O���!�O����-u[��yq�s4�<� "O���!m�N�f	��M��+��2�"OT��C��fi��	GoKZ	[r�'�"��|�K>����;x=mH���	s��d�2���'1ў�O�rȑ	T�)q�l9��җ'$V���'J�j	�al��C kݓp�6L��'�F��!	M��$��Ă�8�Rzyb�'��-rw�X*Ҍ�	D�[�>lƬ��'�T�uO(���X#��/%p�9��'t1��#<}�,h���2���/O�=����'B�a�̧y�(�a�ʣg��<����y���_���ёn�<0��%����y�� �m���/>F+�Y�y�IסCj`[#�U2IȢ�A0�y��Z&�j�8�FR*1n�$��n�yR*�40�}BӍ" ��:�� �y�H�/ն�ˍ:tZdjb�(�y��ޫ+&�Ȫ��N#�|S��y�`ٶf.V�33��.��$���d!�O����=n��A2��-4J���c�OE�@�2lؽE�R��͎#��� ���2O���cB�:�Ձ�n��^H��"O�ŊSfS�+_�݉ Ó	cb�L�d"O�����
+^%���
R��%�P�'�ў"~b��L�Q��}	)

 ւ�RC���yb̟0>%���/M�Ayã����0>	WF��Kh L�ä��&�(����c�<�V��^T�(�!t�@d��h�<ч˓�7��|�b�؅jK����N�<!��V�	H�����5U�l�A
J�<a�kN�t=��a�� Flq2id�h�?ɏ��Obu@�Ɖ��ۅL�7  �"O �2i۔:�yxD�J1c7�|�'(az⩕kz��&�J2[����]�y�nä!�L��C�;�M�cOϴE�!�� "U�F�2UV\�3A2g��q �"O؉Sbc�J�@��]7��t��"O(8�rk�x��J-ٜ~�"u�"O�����@Z؉ �f�"z��H"OJ2 g�*TJFf�f�J|{�"OZMz#�E9	T ⪈�7!�E�P"O�HS*OoP���IƦ6��"O�tK��;h��8�C�4`��V"On@��ƕpf:�b�?VQ��q"Oƀ9����]
��'��@��9��"O���E�b�B(��c�V�b髃"O^�b��J37�~u�s���B�TYS�"Odyڄ�׾?�,��
��h� "O&�{t;xXp��jЭU9����'��'�az����<8�P�$D@�6���$�G��Py�(��C2m�����W@M���m�<1Tn�'9۬@��C�\T,}Q�,�C�<���ǨvitL��� �|i#�Dz�<��(����.�
$�<m*T l�<� H�1R��%���%)R\C��$Љ�3�=`y¯ӫ��B�	��捂�h�H<�i��-M�nY�B�I8)�T���`UP��Z��9!򤝁2T41�#��"��`(��@��!�DF�X�nq��-I! ��˵#7aR!�o��y�DJƆ%���P ��8!�d�*b����K3b��L q�-%!�D��h�L�)5�F.�d�m�*!�*xz�"r�`F����bN�On!���4%�7�. ݘ��_�GF!�&̴QaD�y�AK��<F�!��J� ��V����\�r��zn!���h�jLb��A�$(��}S!�dK�q��o7�N��deW�PX�	w��(�� ����:�@	���
K����"O�]��j[;�<���Dp��Db"O�m)�h���9ò��i����"O�p{eG�)��%�@�P�B��y �"O����ű+��Mqe�H�-�ޥ��"O�`Q�ō]�ݘ/[�B��8��"O��s���6����L�`��"O�TH�.tu�\''�R�X"O��DEӘ:(��e�\]x�CP"O�!ې�ˋ?�U���9R_ԛp"O$��������� �;-H ��O�(q�&��U����%HA�U}H���0D�t7@�;��d+�h�Z,F��).D��Rl��-7��D��U�8���+D�H`��ؕ�  DcQ,k��4!�H)D��)���+S��BM�a�l"!5D���v�P� K��S+S�HQ��6D��g�N�B�q�Iҿx ��;GO44�d`�(G�a�BP	�B[�D�h��OI@�<1��L|���������g�~�<�E��HGąq�*s�La٣OR�<yag�8AbU�'�!x����r�Kz�<%�F��p�u�ޞ<�hL�BGw�<9��4��(��M�'����wiK�<��@Vn�,1�-͂sr�5��I�<qrhJ-S��*`$����%kED�J���O�&̠P*�)H$z�	3憶� D��'w��+�	;/��E�k�Dyh�'�-�p/SE�h Ϙg��Qy�'[2��⋪R�p�AQ��6�A ��� 
�[c�:j}i0��F~B���"O��R�/;C���g�@�__��!"O�`�C*� a�(l*$(�6C��P�"O���kܡ	��tR��*G��!"Op��5��F&��#�B��M��v"O\yy�j%Ybj5�jM
�� �W"O��1�.1�����G*?���0u"O�]���{�f@x�Շ7��rb"Onxrp�SuO�����[�),�B"O��¾h\豉�H�9BF ��E"O�1�e��"��`'Nx0"O�\�FŖ�-DR�qbE;OtS�"O�����ք0H��B���n�"O��� �5I��	��]lޖl�"O�i�$�%;�TPi���^y�鸴"O�����p@��0�����yb�;S�Ĥ�!U�E��e"#�8��O�#~�F��+ .�&��>Q\�#2E�I�<ɣk�6]�갂&a��_�|��G/�n�<ib�ΜS��]BQ�D D�j���^h�<�p��$���# �� ��nK�<�Rd�:&妠y������H�C�<�����t�)uBU�T�8�OF@�<�r�^!r!\�"�(�[`�Q�5����#��'�(y�8۲J��J'��ȓE�(�3cb� }���A%��	dB��wP�dN��}�@�a�lą���`��ł ��Li���&.��ͅȓ�����Z)}���w�;>%��ȓP:Z���%Q�?��9��4 �	��V�����L2p�P�#�.�/z܅�x�z}����+�h�y���Q&�ȓeX���MS
i7�A5"E�le���ȓK3�Y�J�g�zݘ�D�$4��-��C \�؜B����F��Y4�h��@��%�5�7	F����S\L���'
d��AQ���)�g��C��8��1ib���sG�ȉ
�C�I�	��a��"����� >ա�d@�B��)S��9ˑH�?A�!�Ǉe�UZ�Q�	rZ��Cj��!��.�^|�P���DI��P���!�䄩�¥�㔐;=B�Iܚ8�!�oE�1`���WT�T�$h] [��}"��`z��T춑�!��t-��8D��*�ʊ�?��PB���,��!b�:D�L�f֚ cz�
�kZ�4=h��I<D�|`�����8c����~XF�t�,D�Pp����B�J�����3.���L+D�d���P����@��]��ɓ��<D�Xɲ�Gb��I��E8v��5J;D�42�+M9!8�E؉RY�P�3D�`��d�����,2��H`�2D��ʐj�AyL�#0�CRwx����>D��� ��%{f�f��{�)#?D�Ljꏁs=�5(�P���t���(D�XI�C�M(]ra��8{��bV�*D��$����b�@G�d���'D��`%��
X	n4IE�&�n<Y�d$D����!C�{MT) '܉%n�b�"D�xȦ���V�ڭ��I� e@���b5D����J��lO,0�a���.�Jp#�� D������I��0��n^�"*D��#� �7Qr�D�&ExS&Q[��)D�� �}���43 �ӧK�:Fﺵ�P"O)0U�K���t��[I��L�g"Oށp2��;WP9�vɔ�pk��A�"O��RR%UU�T�1��5�8�kw"O��!W�S�/�n����� $�%a"Ot�
R �F#R�i�j9�k�"O~A:cF b'*��Щ��<�b�"O�ܳ��N��/Ɛ#��iE"Oz�RB�I��9bV &��ݚ�"O��	�Ul=)�/�>aG��z�"OVI��J�_P��#�ͣ6����"OH�OIAnV��EL�5����"OdԱt������g�U<:X�P�"O-HP�\.mp�M0��V�J��T@$"Ol�GF��G���b�ϳ.���ip"Oz)�Q��9�Љ'�?��4r'"O���p��I_�aR̀Z��Ұ"O�A��K��Y�hs��]@��Ũd"O
��6dզ_ɸ�Z��~��$	a"O�Ջ��U�eY��FW���k3"OXz�) �$!� /���3"O급��o1�i�qj�
N@t�'"OH��s�K�d����#� H�E 0"O�H�d��--��qwc͗'�v!�"Oڽ�"E��My%�#� �g�$D��XP+����P8Q+��>i�܊�.D���&��8.�M�t3�KҦ+D�XebKN�jU
R�ޒI�d���#D�$"b)�2=�d�&,����P���!D����z����V��0EJb����?D���ЪD�YxFD�5��:�@Հ0D�d;g�Ƣ��� I/`�	Ъ/D�l20)���a�t#�j�M!��9D�� g�T3C�tY@OI�N���1D��q��;B�p��d��f՘����.D�*��U�ԡqv��n�8(�1D�D��DިX"��DBF���� .D�@Ar"�-i)&�7m�t���zą'D�(K���0��p��*Fd���'+D���j��T�D`%d�#":<iD�*D���gx���G�K� @aנ#D� ��i�s�l�)��ّ$�Hi�. D�`����R�Ji���ʦF�Tດ ,D�\���}]�щeȍ��v�r�+D�@����5
�Y���l1�GB*D��X6f�+l�����& T�#D�p�HǙ�H8b%��4�>�pL!D�LJ҄�kj�8�	_�jE�?D��X�Cзk���r���aτ}�T@?D��	�g�*(%���<�z�P���yb+��N�jB�ݰZ��a��y�mעE�&�!d"i�PڤaC-�y"��(�d��ʏ
x�IQd��y"���,x1����/7�r����ybo�i����蘤ĎQZb��5�y�k�R�<c�F�}H�M�A��y�mV'(:\�pL
?�@���ȏ�y�n�!>���qBրiϰ����yb�M�:�@����]�<���yR�S%��0�`�"T�ԱI��ݼ�y���;� ���hO�NNtl���R��y�C�������@���w���y��C�Gn�PD�"cX"'&Y+�y�E�nJ<p)���rYБ��N�y
� V���F��q#�Q��NI�c�(s�"O���5�!b�X`T�\���Ys�"O��"���+U�*�)�b��5�"O��� �Y�4�n�3���,���K�"O^��)	�>!tt�d��"e��"Oْ���T0Ĩ���Ȕ$��q"O l@3�K?H����9w�4��F�s�<iD�#���!��C�B d*�OW�<RK YƒѫRlx���`��~�<�b�S�'b@����uz��c��P{�<!p��jdbyv#@h�H�&Xy�<Y��T�B��i�+P��E0$��r�<Q T�e�ry�Q�C���X��/d�<�lBF��}IT�b�����c�Y�<!��˷��q3��V�(S�KS�<y�B߅E�X���.޻7r��
VFj�<Q���A��P0�V+�m�.]]�<	0.B
D۰i��-K�lv��KU�<����c� �� EkG�]�!�T�<1�g�R4�K�I��ʭ3#�V�<���5#|��s��
u��~�<Ie`�=�>Ɂtg��=�L���C|�<ɤ����0�6��:�݁�z�<��
��e?��A���G.��A�@u�<�e�?/M���O�b"�D���y�<���ʪ�5!��06��uJ�w�<��+��x2�h���y�X��3hs�<AV���$y��b�ÁK���ɂJ�I�<!�"�{��Pw��&�EO@�<���U1L�Rа�$H�7�)W��S�<���%��|Ӱ��4G�h�q�L�e�<�*A�|��z��JHV��d�d�<�Ї_&����h#T���+�b�<�p�ݖ=(��1!.[����Ty�<a)ۂ �@T�V�@46\4�"䀛v�<єN�rGv�R�g����R���z�<u��cLf%7A̹4Q3#+x�<ɧ�ڐ1](�����k�R�"~�<q�CH�Q-[�iD� hU�y�<��"_7K����J�0^�ĳs`�q�<�q$^(C�P]��&,'��VJ�m�<!w	�;=(ҵ	s��q����F�k�<!��Y�䈒`�${��ä`�<)����G|x���#X���s��NU�<�� Zq����'�'9�| ˶
 N�<��,=�.����čF:�b��G�<�j�	(8��]�M�4�j��|�<6���,M�\��8d��)���v�<�E��q��Q�gU6B�t����Io�<��G�5��	��95$<��W�<A�׹�v�P�e�87�f�P��i�<�d��Fܬ���߷������}�<��@�0tn�첐�]4s���sB+�_�<A��ֽa�u#��I�^D$�;N�W�<G�l��)��ލN^�L[��[S�<�F�D�Ŕy#狐�"�Nq:�u�<�'�P�/H<Iu�M�P����q&I�<�d:)��-"��P>)��KJ�y�<�RG�>:+ ��f�Xą�g�x�<� ��O!���3B�<N� $�BAm�<A"�";R&�P�߾(�J��e_�<!G,+���K�ü��@�#��R�<1S�ˮQ�:d�ů$��()��)D��ZC�C~X�Y�С��ҡ3�&D�� %�Tb�!�eB�OZ%��P�"O&@�l�/����&8&�P�0"O�
�k��;�@�t�boma"O�SIW'@l���C�\(d9���"O��r'&���}�'K$K "��"O����3�0�!�ڬp
v�Pp"O�� u��L���j�W��y�"Of��/A3t����nʲ���"O�0ആP�1" �2W���p�`�"O��� @�,"�z�ȁ��'�� "O���Ǐ�7��D��+���[a"O��!�#7�+I
	�^%��IUP�<�6��~\��҉A�൛��PV�<9�j�)S,r������AʘS�<�&㚬w��\����6��P��BO�<����6L��@ຣ��^�_`.���C�Qs@E)b:�)��-8���%�&�s�D�g��Ļ���U B�I;-���8jZ�A��d��Y�9B�I� rx�B�E@
c��R�;��B��N�XL��9qj~�3����2��C�Im&mb���@@X��K�@��B�� ���� �6u�8	�*�g�C��2�)�N � ��� Fڧ^�C�&Z欑8B�_�sB�d)p��&��C�	�}��`����R������)�bC�	�<�b�{G`ҟqd`��2Đ0�8C�	�k�lk�"	�#�j���*C�*�C䉈~��a�t�E4�:=B�BxO�C�I�:�H�c��Eo ]�t�A�0�C�	�%���ru�_e�(��A�b0�C��3 ���΅��A��^p�'������J/G�*d�
>s����'D:�ʁ+q���Q�jd��	�'����/v�tq�ň�f����'�l�ۂ��`��Qڴ!TV#!��'�D*d��`�*��	�G@b��'u6H��@H#%L��`��A�.���'�:��T����F�P�k���'U�U���ŗnGXh�e\�`�:�'�n�ԃZy��(��%���&���'l¹ʗŏ+Sh(��kP�l�ԼQ�'�������5��x�g�7a�(��'!n�Qu	̾zj����K�\�	�'�����9<�(�b�l	1VJ^(8�'� ���бM�r ��L(Hy.I�'a������Z�����l�>F|�Y���d؋�������K�XE*3c�6`6�I�"O�T��kR���Rq� �"O�фKY?x����4,GԱ�1�'�qO�Ȳ0��}�b�r��ۺ^�v��c"O������"�=	�V�"O�yaDÓ����X�}j:&"O��
��E�]���7���K��'�VQ&��*ǫ����X���'>	���%D�X�'�U,Iöq� ,6�E�«'��f����7*�y��=(e�Q���Yh@��d�<	�O���D�	c�ʼ��iώD��}yd�'�ў"~�����tj�����C�x����k���y� �F�1HD�Dr�-s��Υ�yR ��F	�yãm
EKr� ���{�����I�1(����
���eX�d%v��%"O�Mq�)�23�\HU��A	���`�O��Iv8�T�⁏"�j0r,�1��@1�7�O��
�O� �Q�����y�R)�j����Bv"O��C��Ԓ	�ڑZG@J�Yg���@"O`���C��b��crf=�ɓfFPH<A�GL�,y�%�7�ޟ I�m4��̦5�tW��'��ϸ'�ܠ#qiX�^C���3�[�\T@9	��y�DI%�Q��6ݼ�!U�5�y2�=�!K�D	<:1�!�������>)'��<ɒl6�Ve2��̖#CT�R6	N�<a�����уU�Q'n��1
���hO?�	�_��r��<�������wB�"�Iad��d���bJ�6-���(O��%ړ����*фn�����W�ww�ȓT�4���}/���R���i����>W�r��L���(�B:b&�h��o��D����:U) 0�"�E��,l$����	�-L��0䋇�fZ�ze�/6mR��$`�������K��Y�K
؎v�>D�|s3�؊{�x����N/E(td21O�O��=1����4�d�@i_tX1��a��s)�{��dM�Z�(M���y�A�SaX�v�If��H�Eص ^7 ���S�Bz�\��@]�8E{��Уn�2Q"#�͢{y<[�̛+6�!�� �~ċ�L�7
��q��߹m�'*�|be�-5��<�=T^��8��9��?u2O���� j������Ȣ	�s"O���l���.Ы�f��;�"	���Ie�OuH��ҁS��?^9)���N-�S���5����@�-Pr�R��=��B��H�$�����[�4��c�݅��:��/ʓ:��>�i`�:��M�O���t�������Ұ?���H3!�� 3�@�?
"�Mړ�s̓ʈO�OMц͗ ���6%�.�I{��i�ў"}���cL\�9
�>2[re�s�R�$e�G}���*#�� �i�+&�P��cH��`��G{J~��G�/>HPҊ�9QT])�Ri�<i&�Ϩ��&���qG�5Yg�ͥ��d%?�N<����!�$u�a�V�z��U'F(3���i�OɲE��˾�: ���O����<�ߓe.Zd�����:��`�R�bt�%��Zs�)�Ot��2��'��c2Ț�Ln�?a���J�b�שG1qfܨ�A�f!�D�*JО]Ç�]Nκ��G�M�l���w�d+}��iA a��hʶ(�&�@�a��43!��=S���kV*R ׺@�A�U:��O�'��ϸ'E��TI0�-��Hɻ}����Ot��,]n����S�4�b}y��@��$-|O��A�rh��=K�N�#��ǳ���	Fy��|��\�b�~�e��6i��]󥍐,�y K�j�	�%H*b�D�������$�S�O�ؘ���h�Դ�fB�T����y��'R�d���@��i�T�0S�:�'�����)1�A�s�N�I��h@
��ēn�6�y�LV�|�y��R�k��͓�~"��0�'#I�h����*	goI�P��<��'x�O1�T�J�Ú�A�����\��aG�����	�+F^�@��pڜ��V(_�I&���D �I�Eq��[��L(���؅HJ�1��B䉢Fͼ��#d�G��W��%q����dt��nZ3bXe����2V#Z���� 2JnB�I�Sw�Ixc��[�>}��d�5
�8B�	�&���"��HJO�m�a�<[@B�I5O�$�SQ�%-~"�f�E�2�$B䉳h� �q.D-,�(A�rJ:d��B䉮QQt���� 	���+u#�&��B�)� ������]�f�C'ʪ\��IN����*[f�8FǇ7S� [$�*?`�*�O��d�	�NI��s�^+V>L�aO��$�]�B�G�g�P��VL!�{���P> ���6n �-�ZtZ ],��ta�)_W�O������Vo�ͰV�@<�}�}B�~��#�����mO�ej����I����'ў"|�C'5DS��(���-9	���b��i�il�la�����*9~j�c��ʠ�ћ�@=;!�	���H8�`.|�9A�NY�ur�Z~�i
Q���'��zV�t�8��Wi�<��S�'^�Yׅ>R�ژ����<s����d��hYQ?���gZ�,��X�\&����W<D�X#b$ӈr�FihF�D�0&8h#����#F�)ڧ �#p��fS$��+̪a$ZŅ�	hy"�i��2�!��c��-j�,����iX��cVI(m|�ȓؔ*��̡��<}��:�O�(c��E� �0I���ƹq`>X��'�ʓ!�"�[�)^�e��C�ۮXP�d�'��(�Iw�'��t�Te�?�$U;dJ�
h��r�'v�r]SwJ��ë]	cM8`	�'`�yh�!��
a�O�0eў`�� @�$�<r�^([g�[~���7� �Bj(��D�Cmۯ8Ѯȇ�}ƍ��Ҝx �ЇmR5M��݅ȓ#��y`�)�0o�����o;��'��~⢂���p��n�9��x������>�J��iwHɫ\<0��LK�m8��4� D�(
�I�%�acRĆ�o<��S">D�`@V�א<F�9�F��9����h<D�x��ޕn#�����! Լ�G�W������
�@f0�b������%�.b!��̷0�LȢb��.�0j���OL!�!%�L�Z�'�S��8���,�!�d���ehsʓ�Q�bt
S�C�F�!���0;��ІI�R������!�D�?&�t{�E�12�@�!��7v�!�$C�u�60`� �$+ 	ᎏ<�!�Y�WG��R�Ll%.d�EY�q�!�V��B�ۓH��*�+Q9[�!�dY�=�1�W N�G�xu{�
�}�!�$�+�T�7�ЋUG���/M�!�DÓB� �ȅ���{:@|�!
��!� (Ӿ%�!څ%�d�g!���!�ؒkFV(�TG\�+�|y8���<"�!�:S6�M����^ނ�����x�!�D˱F���q�
�(y՘M���!��F6��6hL����SȄ��!��B���L�6�� 2�{@!�$��S�*��P�Ö%�(	����
/!�ݼٞ�k�L\�s�ു�*EnK!򤑈f���jfD�1s&�{��0:R!�䀰�6���Қ��B/�]&!��L|Q���ɾЎ<{��	[�!��'j��4����ܰ�C�;�!�D1�\�h�b�2�vp�֥5�!�䔃V�����iJ�����F.4�!�W� ,Æ�	N��cC�C�F�!�$��}��I��(]��
(#!%�?!�䗫�N�9B(��jBL@��!��)l��{2�ߺz>"�hP@\j7!�69��Yi6+�3#)L�1#��6!�D�� ���U�
 �c����G!�D.na���S1�0s.��u7!�� ��`�]���`/�
Lڸ��t"O���㓕1�ꑪGN� Ϧ�D"O�-�j�0)��L��x�D��3"O�栔�R!��S���>ΐ��"O�5�C@F�d	
 r �
PV4@�"O*�k���(<PafG1Y;NQb2"O��[ώ/�ʌ0bEB?kƔ0p"O���Vo�"*�L��F��Q�^5�1"On�i�-�~��AIV3y�r	�@"O �{VM���C.�o�<A��"O����.�+ <���ң
GCP�"OX<��� ��H�2)����"O$���^I�6TxpV`��l:�"O������k:,��d+W�Y�w"O <�dܸIP� �C�S����5��<T�謉��0>Nر�� �U01Oj"��D�Y�������0�H��"O0���һ��i��!ɳ�"OR�#a��,SIP�v�Їp'�l" "O����G9����Eΰ> ��"O��{��[�$'�����#kY��x�"O.xQ�"D�C{����E�8K��J�"OP�x�Ħ�X�ț)�-��"OZ�0f�E2"�[��� �"O�E���R%�|YTd4����"O�s7�ɾ�̰J��P�$4>9�Q"O�5�Ra�T����I+ �!W"O�!('a����Hsb�G�Pl�#"O�雒I������h�ٺ"OQ�6�_#�B�I��/�6H��"O�t� ��]դ�� @�t�sR"O�0�k��/ݞi ��[�tˈ��"O�m�f���و��Wo�2B���8""O��(�I k�B}��.�(H�00u"OB��C��U:�[�0<n�"O�׏ X�T��,<l#j�*O��{�ɒ?�v�3��Z��i�	�'y���	A7>fPِ��P����'} (���_c�lz��E�8���i�'���eF�9�p@�ãڣ5PFi�
�'�0�#ɜ��5ȳ%:%�0L��'���"���o*���j�&�:\�'�Xܻ���a
��Oe�Vܨ�'�x�&�J>2M�Y��.sȨX�'L&�p�!_ ��$�'�����'�Ii��G�77�!�jD��05��'r~�ۃ���*	�"Q/&�N��'��U��.V%:-`� V&h��'��|���2{tbp�cF�h�Թ�'��xI�T��@P�c��\��5p�'��%��!i�nݰ�"�<R�
���'��'�ť
�,۵�б>��UR�'�vq7o�!H������H�-6�i�'K@�3ŉ�0��Y��G�>���	�'ߦ��T���� �" &O�$�*�"�'�6��NK�-n�}��l�0b��a�'�r����԰w���r薧iq���}�)�G�.�G�T��6T����
-V��V� ��y"�C)k���3��\.+��,���|W6��&�/�$��(��I5U��Ay�'�oV`�7햕3.�C��"Xa]��E�o`~9�`���.DY(֨ ��|�'՗K�u�S
�\���ȡ���0=9FET�s�x����� '`�B0��bM�;�e�5+7D�|	�9%R:ՙ6
E�EE�����1��5GB���3�9Q?�rպP�@�ib��_��F�!�� ����.oH�!�� $�<1b���7���J�pJ�j*�g~�I^����`�x2Q�֊Ŗ�yr�˴!��ف&��+5
�h!뛂We�PKb�m���I;R��p²�C��b�#�=$���̠S�~���g��~Ro�\�#4��F~>�p�G�'�yr%�@X~�a��T!4萀���'즑�P �P�E��T;:�b��p(Q,)�p�� ��;�y�
�fb�l�����z�����K��� F�Lf�d�	
>�Hh���⚩ h�ˇN�	��D��I�̓��''��r�ƐtELљԠ]=[\�aJ�r�4MK 0�=�c�E"�$�z��6Rb�D�]��$��-ԙE�U�'[8,��&��Dbv��%�X2�9�/O��A��:�`����"���2Ƈ�;4J�i�%a!��������B�~x�qT��2e����D�D&���&rD���ޣ"��,��(�����;D��S푞�J��XA�}R���'6�:�Q�w'����c�\�!�D�&1��ܐ�.[~F�)2B@i�旙>ĕ3kOH��s�,l�""�0on:5��&�/�@�$"O*4���=<W� �ce�e9��ٲ^��RDМ,�`4�1�'Bh5���U#6���D�	�w$��u$�`��Ή/e5Ȩ�#!%�brF��,���0�,4�����}��\d�L!QLQ�2�!ғh
\p�uH<^x��?��".!�� 񁈆4L�� R)>D���̈́�cɄ�� ��"t�<ْ`~Ӧ��Ҭ�JDA��N�&Y�G�ܴ5��eHe�
0�9v@�|m���!(�F��U��`�1��zk��j@bj�̝aeJ�kFq���Zi���$��p��Y CȊ$DN\X��[�t��O:p���ޮ��'�<l��n�/z�$�i򃍒���6��
��uʃJ$9�4�'A��>ɗ�'&.>y�4�12�Hc"��~�tdB��3�H�}���DE'����Gj�D A�w�� �G���ع)�pȲp�'�a� @�#A���Q1NZ�k�r���.�>-:�H_��M�6��[�7�@�D��#��	�=X��ZLȂ�!�!t��z���l\�r&��<)e ��P^0���/{	�!�7�.U
�e ŕ>Q&�3����?e�D�3�\�R,�Xg��� <v㞤��Q��5��	�.Ա�!]�R�=:ɞ����C��5�'�"��4ʸFj[�?7�0�R�
"d�Y�H�`I�U>a80�L2W�z䙡U�PX�e��n?vI{�#�r��b)D�\Q���:�4*�&��
�d7��}P����!QlTa�@o�rUdTIH���|��F���K�,P�H�(�#��M�;�z�R,N�A)��D�<�3d�#d��t��-��,�w��=F�1JN>�W�D���d�tp���rMЃ@�$�*��M`�qOv{���1qE�����	�w�T� �A� /�>��e��b� �`�U
a~��Εd+���!@�Yv����a�Ha�By�ɫ�H��	�[ ���ĩ/����O���B��#ky���)�=k@����K*+�~�����л�1�X��E�	=�b5��j�4�̐��"f����M99ߴ�а�� ƖE���9��
z�0,�@	 �0D�,�.
*�]�'�8���гnY&|�W8F�TXBa� 64�A�ȓ=A�\�菾\���5�B�=�6�'~���7���8�D�,v<ڃ7��1��P�'�e�~p�����!��B�ɌKi(�q���Vxt��� C%��(xT��+�=Q��_8L�0�̓F�ҟ��B�A2��E�EM
Y�dE,!�`�`3�ַ)�axB�Ҧ-h�;O�]1wb_�#H����EA�7��R�!8 ä$����?�7�.`��3r*,O(�S���X�xa�%�$J�-QX�����V�/�<)��'�����)[�h�a�R$�d>9�2��!ͨ���Q.P�,R���O��(3��-K)>ѱ��t�� #�ΟԚ��LAr�)�@�4V��x�$�.N.4ٱ�dp	B5�,-�Q�0�P�@��ȾO2e�S�'W&1����҅��0,���⩎����b��WM�][^)/�� �M�dM��x��]**��('��P�j��Bn�lia!��E�	s�'IN"�J�F�	#jIJ N	����+̮2�|�x3��p��� ��I
K���j�֏3���������Lo�~c���`b	)�4�q»p�z�'&� ��GD?��=��m�8��5���LsZ̓�n�]�����* H��q��ʞ�RU��h!P�l�0/PX�;

�,�z"Gסw<2�(�'�j�����Ewtj�cӍsJ�H2��d����n�'�4�]�r��q8S%��:��� T 
6+�$:��u#����8��'��eR@���E�c���)�%�؉���6� �QT#��0��1AB�]}�K�,��C:�yCi'�؍�'�'�
�y���2���B;O�>0d�����̒�xr� 6=�u����r�i����S�Xt����%jn�q��ɸ���Y�FT���G"�001���<	i��`Ȣ`$�G��'+B4��ӡXf���'۹,wbyr"Ţn����.h���'�")H,�f-S [n���V��8,utY*�w��	;2G^@�z���o¹��0��"v��`4)��=�(��	�`@>L�5e��$�\:���79,<�KT(C�[]6I3��wwz\�3B�=E�:t���5'�X�]�����4/�"	du�B���H�P��-˛[L�[���\X�4�f�Z0���!��is��U�5(�$����Z�rPY����:h"i��B�[K��ᇔ�lsԔ��&R6.�0���D�>��f��1��Y�F�U8h��!
��*&DC؍��
Qd��2D,6M�#t��A��AJ���(֣ɆQ�M�B5YM
�[�+9q��H�ȍ8z6d�5Dq�p�(�O�`�Ç�7\D�s�K'�I�_��1A��� $\8��@�z�ꍻ務Ӧ�2��
u��i��Y?v�dB�B�GE�DP�.�����C���*Y�T/|���C��9+$R��Jw���7M+?f
��,cP� g�4�]����r�E�s��Q8����DJ��YA�N-`V�����u��P�rwJ����?\�� �صV��LÏG�pf�:��'��\+�/G�qg�fU.��̸AF�F��<�q�I)ybvA���	�kp�Adi�2����V�R���1�F���X�&�V4eS�� ◝ ���X��+�ɝ!���H�0OhUc��I�(r�Zw8�$�)�^�0��`'KC�yB��W���"��
MU�T��E��{"��
YX%j ͈�1�C���򄁴!��,2s�ɖ�M�	E�/��֤Ch�=�҇���R3����i�C �|=�I�2�w�<�C�I�%���Ҍz��xP&.E��y"�Q-�"��GKLc�T���#Y^�D���ε8�w���j1+���Ha�=-i�I��'�l�	�I�>[�
�c�*�c����H�5������>v�6��	�y���	�~�?)Q�_�z�D�i��I�?`�����J؟�@"�Gm`�j`�N�0�^�f�]1byx����.P�*c��`8�X��,u�r�K�+7ޞ����+�ef�K�##j�R��ƬE=��df�*^(�0�ʨ+(�T`���y�!��K��P��ϞA�J��+���>zfQ���;:��p@���\'q(B!t�ԋ/Z�ɴoռ49!�d�8Y���0 B4r/�-y��!2-Ё���>Q�,[�Cg\�>�OD�p&��9}*ru B8�&]J�O&l�P`G1o�&�j�"ܖK�:@
�t��VK.L��MЄ(��!��8�d�ȓ7PV����֌m-@`��W���ȓԙX���"G�E��R�66��ȓIfh��ַh��<��k�7oexU��6��Q"m޲|��2b�,U�ܼ��l+LQt';h��1կ ɨ<��<�da���e�X8�@�������j�<�"gkT�� -r�U�~H��CФH3�E�x�8E ���|��q�ȓk �|hC^oN 4 G�ksfH��'�Hؓ*O���i�v� ���A�'�l[G%ūRj���4{@e��'�⼩V��n�h�pM
����
�'���Y�
Pi�-���Y�
!֠Y�'���c����H�K�F^�*�'���б�Q$5��ə�f�z���'M����/��]�@)׵r׶$x	�'�
D�C/�;
ZD�w˟n+l}��'EL芕���a��p�L;c�j��'q|�X�H�U2�D	U�#Q�8�K�'L^���!��oi�̚�B�0wb42�'|`����#�|�� ̤-|�d�
�'R�j6�Y�L%�W�������'���	�nEy��@�m��c�'Ό�JlG�"�yF�>pҔ=Q�'�N�3E�ښB ���_,]a�� �'�ث��_�;�H�d���T;PUZ�'"��+�cPLEl p4�xH(�a
�'	��ˑO�dÎu��%��'�xDѠ�Y[�ڴx��?XGR���'�Y)Չ� )7f!#��W��I��'Ҙ��1m�Q8����&E$5������� �в�f�r�\P���ް� 1:&"O*��r RC���k�*Ǆ;8 "O&5����S8��RC[00Z���"O@���\K��T�]���y��"O���X�p(p�BT4|TR���"OX��5c�L�V����'��1�"O�P�fE�y���zŀ�M�J੐"O�@4"�?i��b3�#�6��`"O�$��k܅)����$EU	T�Xm�G"OqҢ�A� ��=ᔯV��͠"OD��M�����*s�ȟg�b�"�"O���g�^}>Ias��j��""O���<FL�4#�kq�nA�7"O�p��/&�Hs�*]�1�f���"O���e��:U���)�{[x࠷"O���3�W)�y;!%���Lb�"Oҵ
E/�n��HYf�^�D�  �"O�i:�I�0F\`��B#յ=�F4a�"O�}�3^�/�n��tlJ&b4�91�"O�!��
mX|U�Č1m=��s�"OR�j��Cb\T�K7E?�X �"O�|�AJ�EL �k.L�e8�"O�T�Q��#-��ep�۠_t�""O~=�[h���LJ�O�X�{b�<e9!�d_�x&*iA����'8P��UKZ�|!���,H�$�T0\�"�h��H�!�$��*�}���)n���j���M�!��&�&hk4�[���x�2ƹ,�!�DUpܰ�Kb�u,��S�1	R!�ĕ$W7΁��t�\���V�|Z!�H�l�`�Ҭհ<�&�c�A6k!�ҢI������\)3�)��iE�	u!��H�2�X�At+�/���n�=v!�56� �k���IVN�	"&V�}|!��ڶ�`T��"H�t�E�.d!�d�$t�F��F��wiT�Yp
.Hm!�čO �łV�Rm�(�ZR�;Z!�,@��� �C)u�\�i��<_�!�ā�:��z��ܩ\6�qu�D�Lc!�\�J�bi�����q񗋙 o!��-R��|�0F�N	,�#��+�!���-���4��E�������?R�!�d�68@��0��U��+��(]�!�B8>���p���۠�q�膾�!�䐕\Nh
��*���E%�!�$æw��G���HgN@�w����!���'�J��w$�:fHq&*�_T!���$+?�xR��\�Z
�@��ȷ,�!���0�3�06֨x�膴F�!���&��]� ��Se��\<	�!򄄖
��i��SQ�g%ѕSf!�D�Z.��b�z�M!CdT]�!��>&ȴB�@� �J�#I!�K�%��S��+}��Cjw�!�à����CH��(H4�!���~�v�1E�#l�Z�����}�!� �4���aDP�G.�3d�)n)!�\w���%�+Vʥ�Ĥ��PyB�02����ԫF}~���C�	�y�8���V	\�~]��
AHE��T#�	�`.�'"�����I͞]"������sk"O�l���R�}1�tC�ӮW)�E6D��/(�$�@v�<�B��� �SFpR4#q��U�<	�&�F�s�I/��ʒ� ��y
ыĹu���� �3�k��=��)�!��D�q$�'�Ό��-�
Y$�0�O��3V�֒���0��*~l����\�00@F�U� ��rX&T��<aS��$yX� ��M#�'�u��E�� 2�0B͡?��q��)s�T���B{�*,(4�X�dXĽ��g�7Z(�'˺�+��D����94-�+���$I�s��6D��*RF�%씈��0uA�Df��/ b !9H9iS�|�M8y�8�Q�cҌZb�	��0=���]�f^	�į��K2FLU�Pp3m���nL�(7D��
���=�v���N�`�����2��0g���"��+2(Q?��`��6R^��ՠ� t�j0D�{T�X�d2صy�O���Aq��B��}j�>�v"Ba������Ҕ�P�� m&��u-�<s!��@�/��Y��ص��|�&	^x��2K���,����jqO����h!���KF��,g�@��Q�'�A�bk�;~�I�Ho
DK��M��G�:�v�<-@���0=a7�P%�� �%"�e��l��Bl�&٬}�0�=�I�-l����;�B(A'�1�܌��GC�{ǤY�Ɠj2��@Bېc/�	Yd�ɸ*�-Gz��4l~J��Hq�'(�9��	'�H�c�,q羅�ȓ5�XR@R>(t�Us#��+�v�n�I�x���O?hl�S��M�9`>�����+�}��PB�<�QCTc��@
���4q~�U�t�Wy}��!@0�����dx���p�ށ
�%㒊ٮuhƙr��:�OԘE���0`�;%%ݮfa,4r���w�^�;G�Д��x�N����j��_ZK�h�V��
�HORta��D�D!����#��*)Дz����ʞq��-�=�yR�ȽKX ��3��^��S�T��ٴz��h�1�',�6)!��
y5�?7M�z�؋�D��G�v�ȕ�['m\!�G�0��uڗ����];![�`�p *��Z�|P]�gJܷp�+.�����1�_�POR����*3�8!��<�I�"fZ�SU�d�!bP�{%��?Y<8+�Y�a���e�L�h�<�C29��	�'e�ts�h�'JIj�k�$g�����5�by&��	p�l���d��,d4d�ۄ�Ֆ5 �N�t@�'XEL�)���>\!�$B�#�֠d_�^P�}3����"�(��M�3D���5�6&U&�a���ʦ�yW�H?��b>-���]z�ae������r0\O\II�@ mm���'��IWkשKRH��&h���D� �q+7}R����@"�[��@2.�2��V���0���=� 'ך�V-*��?�'��I3Dj�k�@%�Ba\/@���o6E�N9��L4�OF	h�*�	!��a��P g>6�� .�q�F�82�>!u�|�ϋ,*���ɴ>�_E�8ɐ1��{;<Ћv�ƞIr!�	�5nxi�p� 5)L��E� O�xr�Ɩ�|y���r\z����g�d%���h�#"�E1؈q�D(�T��Q�>v4r��"�y��+Z��[)p�x`A+3]0����|RL����I3�XY��@�]���s�̜f��<C6�2X���xw��6.J��v�Dƴ�J��Z���l�$)a<��Ĕ�4�^�IF��H X��#�7�DM`3kU��7Ñ>�P
�Y��2H����q�޽y����v����9�l �Pf\���I�K�|�s��'k��R	زW9$�3�B8An��	�'
���!d�1t�].]#	�'t��FJ����`!*E� )�D���$�)l�2�Z+O�L����lJ�t��"'�,���0#�h!
�'y��R�B�.M�� �.�lk�Ova��Y�j���	2�^����g��w�D��G�%�4s�+�����s�X�#�$� q����Pf�<�E��:c���h��ҦHx=0�O�\*�Ŀ?YZ���i��P���%8&I,��s�M�W4���'-��%iBIo�,���U"���$�I�uf��r��i�Rs'H:M02��*.}N@a�foX�8{�j�4?fZ���N̯|P^1�T%�<a��޻2��YQ���O����M��P#���V	2}�%l�)zS^����ic���k�-E�*�e�%$�8.?k�@qC�YTY���������5�U9u�ھF>I�j�Yg�p!3a�T[���A�'��AV����EI�:@DI�E$�3Q��R��S�`B��!�1���L:�$SD�#!j	" ��>�Nd�dc��G�2V�?9��N�V�I%k @�&5`t���`�C���?1���&���!��O
�҉� �� �{ �i@f�v�%O,@�Y"#�f���F!h=�x���؟�[0�OBn�>qǁ�W&6q�#����Dx�*�Ly�EO�[w$lScA���a�.UN[�����OZ��B#��P�S@�[?`�~�3L �T8�HpBCE��}�G�.y�����'jI��ݮGR�<�)Bju)�&�U8��jdŊ�o�*���W��uG�Ut�M��m�$�(� �bmQEbG�ny�� �5eh��B1����<�ՠδgm��J�\&�II4�r�NQx�^��\I��(�䐠	�F/�����x�<0�N��u�@Ah�"ޜ�?���~ʒF�&���1,A=�ּ�E�@F�	�{p�A7K�X�$'�5�w�O�������
�FM�Ql�',�H��Ve[Z�T�{��T��.M��kԺ��As��~�C2	�Z���Iӻ~�,a�U)�v2�9��=O6�����^�"�9�㘳
�T���is>i���y��#ڈ����8��1��!�"�?1�mȩ/?Dp�#�]�ذ<q4��<fn�ꄜ`�`4���l�f��_(عz�'�M�Q8��@�MS��9R%�$�0����� p��ǧX�B�R�A���H�a!,OZ��#H֢
��4F��v��3&��",ߗ9`�:�"��)�%�G�ɀ*��U�Æ .q/�hʢKаx,��*O��������*$l2����Ns��#��x�4Y����7�I����g	uN�x���S�y��f�*�(���I	�i. �irɟ�>ܑ��KB�>����BBXyR�o��~�N/E�r/�GG���1ူ=�T�r��iB�yP5h	�3 4@6�])[��SuD��|�A��dq�p1��;�ƚ~bqa%'�#DP��Am��wf����<	7�חl�(S��.�T�G��B6zm�v!A
4�L���`$~���{Wo� s�e�9�3ɟ2q��Ѕ�i���"Gj��)�ܘp/H$g�v��	�)�Ԍ+ �Ȥ�?�q��,ty��j��HX0��9W�]T<J��P��,e�$�%�]pR�i�4,O�(���л\�$����ٙb�dAQ��Y�c�`IY�'l���Ý[y����YR\�b�
E�2DS�Ď$���$":ٰ5Y�' 8Qa��n�.dJ���V���>	H�4	��ۙ�?�d�ً2�#|���d�5(P�'HT�
��@K�<��-��&�W�È^�
=��n��^�)���L�g�M�Nx�R��0�@Uc�~B�	��Ra0�c�+R΢}�gC�/\�x�&b�=!�$�"��e�%n�f�&�3P���=&!�$��#	��Q7��A��ё#�]�$!�D� #��#�� k�� J��I��!�䋐A@�q(2���q�޸����!�Q@���ɒz �P4�.�!�ʚg�m�u�]NdYhAM�o�!�A&e��� � '@/�Tr�m� E�!�>L1��'K�x)�&+ g�!��b�ƹh�X<0ab���r�!�DT�J���@D��4u��$��նX!�ƈ1���ҫ�0!�rQe�]L!�D�2IS��#�Zrܵ���>:!�Ė�7m �Ȓ%�-6~X ��J!�dK�&���P�!�; D�4A���C�!򄑬Z* �����:5ƌ��-6^:!�6d�bxb`㚛�]a��ժ%!��;b�db��;f�����7R�!��S>z��H�m��n8���pq!�«{����w�M�ph�fdP�Yf!�d6Sg�=9��ȗ|3�!k�$�^s!�ּ?C��23�(-�B�w!���>(&�SE�M�cz0a��cQ!���/1V�ڇ��\m��4�ȡL!!���)N����؈_f��w�H�8!�$�;v� �@ޚ8Xl����X!��e��s�ϕ�B��E���^�@_!�U�C�j����O�v�<0���A"A�!�h$2����h��Z�&�+!���?)=+OK�z�jA�G��&!��aTp�{sʞ�g�:8B&o!��cx�\)�㖮�dY���*^P!�DM3��u�/)�f���Ϯ@e!�I�j�8�Ç�ЛA֔�j���B5!�$¨s�� B�L��C��L��ES�U!��މ4��qd֌I�,1�UC�!�Dv�)�UNJ-����L2!�Ą�ajnͳb�w���3��D4n�!�� <������tRB�Q�T3"OP�Kd��3�P`0#͒�i�T�k�"O
���ļ/���%ؐ|�ѰP"OPeS��-��<9�N1.�(�Ca"O��"0)�;=���2��(
o��;d"O���D��_V�	I���3+svy�"Ov ���ܣX���ꆉ�.�F�p�"O���'�m��M��ɠcF�s�"O:�����5�T�`�9e�Lң"O�遵���U%pI�@(��/GbMz�"O��+"K�"o	Fp �Z�=5d�{c"O	P��N(i�t@�@�W[n�F"Ox;Q`]�ڼXfТ.C��I�"O�a8#�ǝ~u,,+�$��S�� *�"O\1bD�׻9�}�gd� V�Qɐ"O�Kf�;߂��q��5pLHa@�"OF ��bǪ]Lt�y0BX+-���"O8YKS���3W�	�4bV��	B$"O���ę�xT����3>$��"O�0�d(�?��B"���3���f"ODL�2#L��Hh�\�FP*���"Oȕ��$۴:�d�R*����"OX�ʵ͚�G� b��Z=�rp+#�d��:�lLS�l�/[Բ��`ɡQ�1O>43��J�x��͓�-߫rي9RA"O��p��=>�5(���	�R��g"O&eas�ǜ#n@���F^�)��"OJ�ї�}�:=�V@�2lj:��V"Oj�A���{B*!zeL�-bH���"O��RK�B�m1$%�2Qde�3"O�����1*�v��dasd��K�"O𠺖��
��ʓ�^�I�1� "O�(p���$��iw��H��L �"O��R�o%KɖXZ�A�BO�=�y�@�3-g���G:@����r>�y�L�6_��bG3#ƶ��QɃ�y�똨B���i���R%L�;�+�4�y�/�`�]��N�TXd�am�.�y�?$�r�j�/ўL���o�+�y�	�S����ůD.���$KӇ�y"�ΆdY�B\78�jd�%��$�y�'��.]̓��(Y'�8zb��,Z��a���'u*���&�)�'.��q�@�f�D��Ó�b�6�#rI��"�A���~d�wA�3}J?͢���+m_LD�)oָ\�A��-��Qڤa��PL>���,h�H!�1K9�IQ�%?�� a�z̳J>E��� 1r�a*"j�x)Hp)2$ ��y��V�P$�qd3o\xȪ�!���y��Y3l����a���� �]#�yU��B8�v�Z"��+�P�yB�V�L @  �