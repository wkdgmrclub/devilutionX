MPQ    O�    h�  h                                                                                 �;I=�]
��c�D�	n��K�]�HCpkn��r�HLC.�$2��J7�0;,���f��7V�e(ΔA�6��}O�x�G���W-����D"�j�8��"Fi~���">j�\�w�q��w7yKk�Ҿ��@�NW�� 0Λ�<i���M�3�[-��%���:I̵dK3�~=|����V?�ˀ�v�B�Mdq^��Ǿ�,ҩ�<\�E� 3�ޛxM�}����r�Ȯ��]/�5{�Aq�������(��$E���g�q\	i����6�^���<%I���(x�斷�t$�}�������JUN���b�JƠ�_��5A�S���&\y� �+����ak�I\A�5�cq�Q6�Z�H��!.X鿋	�w���Yq�E샌�h@~W�L+���-�*���"3�I^��]X+���cl3�ŲL����{�j��C�C�!�`Yп;�~3#^xʡE{��ɗzsOr�1v�<�#}�@�D�/����G%e�'D�X�B�T�q6Q���{�u�I;�︝��P��7�	y-���b��f���M(�����|�oq��'Ds�	����ˀ�\���qCe R;ݱ���W�~�v^���5o�o��)u��L�B����$�����>ɾ=U�Q�v�v�zk���\'Gp����jᗳ4t{/��B�߫�*=������W�#���[��]Ǖ#��r/&�mw&M�o`v6&\_(��=N�䊟�A�ì��,/$R�7��-<�wm���u湴�.L3!�ȹj۷��-��p�q��/]�ق���W��m�v�}����r�%y{8���4�����G�y��u�4�n꾽*U�lY�����������٩�$��ڠt�/����ZLqe]1���Z,*k�Ԓ�E.��c�g�A�.�.�~��,՗�{=��Y���Q���sz�tF��ִ�1]X�Ϝ���\i�*��-Tx7�g���3�C=QA��282vnY�N�;�A�s���_���AU�3�S߯x1cW)n�]K���~ݾ�^��	Ŭ���_Ձ�A;h�ԊxWP�=?V؝�lM�?��U�
�-F���u���BK5c���u��1h�j�e+�}�	H���|�#hƓ�S���Iᬐz�QV7��Zx�1�bf8(�U<A�u���P��(\��!�g{Q\ͥ����i�#�΅����ݔA+�;�8�4���u��ꩅ�1����`S�Wk��&)�ǄB�� ����v�3M��<�\�g�����!��ui�� }�+��HGB]"�pUiul ����5�)�s��'�u9��q[b)�����/H�����s�	ah\*�IؒrǴ��%�U�p�1?>!ܒ�Q5μ��}��f"^���\5s�oH��6D���,@�&oω����g~�:Һ�i�(�������^=,4�}X���pN��;�u���$j_{�i��Ue�Ms����|�̺ 5q�拋���i+J1a=锃���V�Y����A�U7�Ͷ��.�\y��s\ĈpGwH8���M����s&B��D~��-�h<K�*S�"���,����a���?cR!A8�)9�7�[F��.����;Tj�䙷 `oX}�Q ���a�`k��O�|ԭ��%ܕ���K[��V����0#G)�[ЫY����4�����;,��M��13�N�����[bG�sY�G��)��x��e8n�'����A���w��+����.��P�lJG��C�3�=��X���K��ҹ:��i'��Ln	���a��ť��?gg���Į�3_�)�yDe�a��];��K�w�J-�v��m5������D�Fm���T�&|G���/�Ɏ�z���^�"h�r����+��?9���}R�~�lAj�m���'�5d�­��VO?�"��A���Dx��o,(�	hE A�X�iAT�e��6������!�B�@�rJoo�yf���+�O��wDac/����EPV�����$'�<z�����e�����*;�������0���,7����y�nPq�����&'ff�"P��Q��?���|������W���kP���B��Q*]/���6R\����=<��[]����� ���@8z^c�s�שQ-�nI|�xk�z>�۲�8q)��ǝp6��>a%I���v�p�p8_I�+�M(5�Hl׫o*�$f�h�ď&3�3�k�	Ͳ�����o܌�_K�9)r��!\S#C�j����)��+1�$�W]��9�WO��XH'��7��	�W������,�V�>�R��S�
kn�Cq���S����R��[�#�V�(��C�{}�h�gO�"k3�>؅w���/�[Vg���0�� b�mtm����Z�Ǉq�8ډj,�ް��ñ���s_�+}�]"�s&C���!g����3L��g~��MT��#W�Z.OJ�+9���[�|xƩ�����
��EC:����_`BֲS�s��ݝ�Jw��G��T�mU�ʙh?)�dIt��<�py��+,�Z�%��&�Z,Q�~�Y'��߲����Tȁ���ݽ���^b漕J�7WA��%uL��<�u3���;e�R7B-f�@�1<�Y�f$_��\́+Q��U"�v�uP2=WVa�G���X�4T����4, `��B�ݗ^xs��/lm΂,V�6b��ܞ?gM�(4k��B�Xg�'������l���zaB2FY3�F{X�NO��
VG�9�:1�>B⏾�dqJ{�����L�o��;��EZ���\��:ᣑv%C�%��JC�o*{f������қ��M9�[�k�9��E1C"2Sc�&����v��=2���gPd�I����X �QGҎo������kN�$!NJ�<�Z�T*
S|Ή��I=Ⱦ��Ĵ$3ŉ4L	[�+v��"B�����]樇�]O?�mu!�֜�W�0k����}5���@r���3꼶�&w���"�Q��+�5j���*��0R�#j�^�a�N"�z���֘uȒ�K����|_{O������U����4�e�VU����-Clo�Tn¶���Kí��������ezm�x�%�t������E�ع��.۳>��]j	�����7J��5|rѭ�;dO���XZO�;�-O!��٤�G��뚸m>��G��MQ�����b�=cl�P�>L[��	ǅ��Sȑ�(���+���~BJjPqY�B!�#��ܩ�y�<׵P�ۓ^���b}����Z/r���->�]��{�M��#Y�T)�(�\�$�ݓkeqwM�i
V���^*.'�I��k���s���(��N�g)�fyw��K݈:KUI���-:JԈ?�z�'5��SrC�a��L<{ �η�.̨k�Z�IaAJ��cLS�6�ŗ�㠇!)�`��6wcm�Y�ū���h�� W�
�1�-���l!z"�W�^�x����+]�Fc��W�M=��������CG2�!�&��Y;�7�^2Z�<�����p�հO-%�1�vĞQG@��(/��"�����ܧ����Ș6,��y��P��;����VĮ�X\�d}��2��}6���_$�*�@���8��3o��2'���	��S�F6�7"��qOe�Y�ݬ��h�9qE���y6'�J��K4�ugiH�=�*��u�B��:(��9���,\B���bzd����G�L0��?t��ut��������=\������WY���k����{��� �M@�먣M��`q]H\�.K������ᡙmNÇ̕�gf$RwV��(.�Ҟ'׺�U��ՉL���Ȕ�÷�#%W�l�/������Ҿr�#m����X�>��X%�m�8�*4q���^Á��y�����n%.*��Y����h{���"��^�$nF٠O7��
*��4eXO��Z���2�E��?ckz��|!������0�#{��|Y�9�Qq�]sUa�F�qqU�1X���Bև���i!r�5g�xq�g(�����>=L�Rߍu$210�ntY�ɐ;�UQs�_���	��<RR����S�d�1~��)�l�Kȵ��w(���.	����*_���AV�����P��?N�靯�H�O�5�
�޴F�G��'�$�KpS�3-/����ő+Dӓ	c�i-�#C�.��WԲ�lV�	=��7��^�����a�(���|��u�z]�K'G������U2�4t� ����c#���t�A���V���(��$�O�@����j��l�>�#}�[*�Wl!������g@��k" �g��,M��R�WM�g
���>.��2��XH������9�]�apP�Xl{�jۯ;��D]9��_��P��Rnyb�[���N/�+���s�$�l\�H��m�}��%� �k�?��8������}�]�A:���5H�u�DbPݳqel�A������.~@��:m��i۶h�=	��Sk�yxO4���X�|�5������u�v0��jb?���"U��`s����Sgv� 0L�Q�;�iF[ea�K�~�(V6��A�O��(�L��N%y��H��8�KpKw���Ջ~�M��B�ΊB��~9�-03�K�DZ�]8���������GJ�c�TAS�q9`M�[!�.4R��ֻ3{?��w�!o��Q;���`FO�������%׻��u�c:�V��S���#"D�["n�0��/��F�Y;��{h��(�3��-:���g�VE�ΔrGE��)�<j��چ8IPY'7bh��T��
E�$����l.��������|_�3��.��l}��	 �Md�����{���E<�>�G�`� �:��g-�q��r�����T�����i]�h$�F��w�1��1v��_b�OY���.�d�m�N�O��|\Y�벍Tɩ�o��>��9�)�]+6r1��&	/?�ٙ��eٙ�ul��f�{�
��5�b���O�Y�˕��\r���f�JJ��D�,E�ADX�}�Ts^�ä5��֕i�O�ֻ��%�{��J
�zyE����
n���aD�Gr��f���?�0���֚�'a��zm���9��e7�Q��I�ە$��0��,�����]y�q!ӓ��f��"�Qг�y~��\�ቫ>�m��������hi�]*��/��R�ڎ�+=�[8���ń��.�;R���s��QH�;I�:�k�E�>����^�)Bx��0
���a@�Y�3`p��Z_�ɜ����5�����>*��f�,?��3�T�k�E��M�����/��&K���)���!׏�Cu6�����,&3��C@W�9�[^�k��H�7:���'��)��(��N> B��Ί[F�VC��b���:��zn��4#�_��N���HX[��B�٪��
�9;KwN</�i �E����D =����?mC���U�ч����Dz����fw���a�d�}���n-�]0���D��.��ѮJ��BL4ƈݒ����U�O��(�V��.�|�v�1/�Ej�E�^ѽɋ7_���������F�sk��3tUHQth:��d�;��ʁ���D����5�Ϟ�ИZ���y��'D�x�mm����OTC���Wʿ�Y��BϕE��7�0���O��o�u�Yz�;Oˍ�p-�	@><�"0�!���yԁ���0��v,A�2؉�a����-��D晠�(,�k����NY�e�m�����tb��#2M^Nk����H�����J��S�a]EY�u!{3��N���
�	9�!&יt�yu/qeЗ��f�x�:oO�x�֕EU�+締:��Cv@��%��Ct�]{��J݊>��y�U�[��9�0�1���S>�]&����:����P�lg�AI2$��b��X�BuG��O4��B������NeV��+�/R^S��b�[�:ȹhj���3�hOs�	�6�+Q���]p	�:�.�X��&c?�A!"Ĵ�k0F	��:�}�@y���ۗ����w&���՝������+�y7�4`���o��~���\��oz���l�����G�k�7���_֘1G���a��J������3cUYSS�(�o��t�q����B8�m�%˼�c��ez�x���t����je�`�t��Fێ��Q�j�{����17�������{�d����3�t�v)�-�$����G#�3�s�� �E	ã�ݭ�(�=���P��Lt{����R���:�M/Գ��ӆ�d!B�"EqT��|>)Ǣg���r<R�����T�g���}��Rыr}ۮH�2]%�n{jyͳ^ ��(���$����&��q��mi�=^�왟^e�g.[I���Z�o�\&������[E�A��:l��#��UDݑ��1GJ�k�� G5SMI���|��� ͑f���/k��I7��AŦ�c'+o6��)�~�S!$T��A��wfY����y�	h�%3W(�|�̹�-MU�Ǚx"��`^�ss���+8�/c��f��M���<� ��CAQ!��;j��&�������T�0vO辀1�G�F0@o,0/��}���{ѧ�z���6G����+��;0�.����������|�h����\�$��;�>!��8l(��o'*'���	�����]����e6�ݧ�]����6��8߽�V��%��_�u��8�p�fOx��Dg�U��ɴ�E�7~�� z�aU����G&D����9�tq|{�-��!�=�]4��v�W��ª&R��������(q����M��`l��\Urˇ ���k���b�N����R��#@�-�P�uO����LL)0��oX��/o� $�gr�/k&�`�Ⱦ���m��3-��I-2%<��8���4�Jȣ�����y|���̓n`��*��Y�xt�;;��_�n�4�$龣�*��E�O��eS��z�Z�[�
��E$]�cF�ᛷ�Q�dR� ��{��Y��pQ���s0?<F&.��1S�]�R���Q�Pi<������x��{gc@��i�q=G_�����2�y�n��JD5�;a�{s-'Օ���7���QfSU9L1�])d\9K����1�ڔ�C	���q��_K!�Aq��ԀͥP��V?���J}�C���_4�
>�`Fq�k�x�YK�������'� �+�Hp	~���#f��2�%�xᢜs��p7M�����X}"(�Ki��wu3(��F�y��<$���7�͛6 뮵�#1�������ac����j���kR��K�Χ�!�� R�V!wW���WJ���@�8h� f������M$���Rge�(��Z�M�T�ӏ���5��Kr]Xo5pKc�l���j��_�����+�z����b_ �5}/����h<��?u\ &�H��*��%PA�f��?�Ւc�J��}D��r�T5��jH�c�D���,���\/��t���f~{:�Ki�o�=ݿ�7����z4O��3T�p�:�� u��z��Sj�Ч���U[�s_'��AR� +���#�����ia��a3rM�YduVq���)�A�iW߃IΗ���y��{�&�?w��$�&0LM���)BO��~T��-�dK�~q�����b�������,c�6�An�a9ۂ�[���.o�C�qC�v�B�Ҵ#oΨ�QVn��B&`!��Os�7��%�"������-Vh�s#�~,[F����lG�*
̡C;���Tw�>�3���u9*�2�h�Q�^�)��G O )�ڃ�<�8$�R'r��P����ʟ��Z1�.���b���W��3�_��<���{�������B�B=�Z��ނ�#�����5��g���:^�8џ�o/HF��V�]q��A�^w69���h1��U����Ӻkv�<~m���J�|���mb��$-������r�+�!�p?�6�{n0ٴ�l7)��As��E�y5�@���}O�᧢�)y�w}��:5*�%����E6b�X�T���_T����c�׈�����J�fkyD�^r����9��DWL�\�!��NF�љ��d'��Tz(��T��e�o���ٻM�D�J]0���,�?H�YF5y&�gq������Jf�7{"�V�Q0���ݘ�����F��u�9.����]%A��+�Rҥx�9��=2��[#=�O�V6��s[yXQcP�Ir�Uku0�>
H!�nlA)T�S^q�Za[�&����p�|_���Do5�@��a��*��cf&����N3���k�7�荥��S,�B��Ke�Q)��!R��CP"y@ur�_@�!U��ڤ�WәH9����ZHݧ�7M�ܕ����l��@�y>f�>Q)�I}8!��C�oF�����2&�y��#w>����9��3Hz�}W��Xj��4��wi0�/=���*;�&�u ��z�mނ��P8��'�8���+_���J��R���}2	��i8��hq�����IF~�)i��:(�Æ�Y���P�O L��%��I��|nyn�Z�4��E7����:�_?/��*���h���b�N�>���NU���h5�Zd�ƱӲ�ϱ�QO�!�s��i��pZb {�t5�'����(ݠ��-6T���Х��&/���y�@�7@犛J��)�$u)�i����-�|�@	�<N]G������!�T��lvg,�2sܚa�s��E�ӷ�U����,�p���z��D�� ��m�D��3bu�y�>E�M��tk�\���I�]/f�#���A�axlY)7({ȨN�Җ
�Nh9�(W���ŏ4'�q���v�h�Sd~o��/�q��EP|��.:W��v[�%�?CO݀{����%�,�ȵ���d[H��9���19G9S��&+&,��펯�:�g���IM�n�ݠX���GH�ɥ�s��J��!S;A�zN����Pd�
�S�4���~ȴf��j`�3�v�j�	Q�+,����w�մf�SX"�j�?`5!"��M::0!�x�r}k�N�Ha�8�2�Y&�=������*Y+޸��KN������}Ԫ���p(�G��4�������_1��=���k��V��R��ۭcU�c�# oW]{�,���Y5���˗'6t�e��jx���tP]�%��{����)�iꮌ j?���B7 ������h�dE���z�ϱ�-����0�G~�ۚ.�/�� ��� �j(��c��=�'2P�#LLϻǻ>������U�����XB��QqOtvש��]>ީе<�x븑�Q��pm.�}�K��g�r8f��cP�]�e}{Eų���f�f�(�@�$Vz���Nq�5�i E3�ǐ^����)*I�kT絍k�����]����huIaݾ#U?����H�JJn醰Z5���S(��״L��\ �t���0�kKV�IR˖A@��c#v66��6�!俜��w�~�Y�0���h�ȵWc�S�gZ-���"2�"d�^��xx+3�c�	Ń~���W��{w�C�o|!����P;E	��::�r�x���t��m�O�x�1�8iĔZe@J�/Y���L�U"�i����1�6b���o:�47;kX���Ӱ���@7�B���"�ה���]�yV��H��l�o���'u#�	�=��<��KuW�e��ݢ<;�|ү��՛�o��� 1���8u��ǈ3������"�p�/����1*�'wEz<멒o@G���N��t�R���\�\O�=���~'W���ع�3�w'T��b�\�M��`gA\p�Y�Br�5>��&9�=�ז�4�R��r��aZ�0��xL��P�J�d�j��[ʱ�bo%/nM��¾��m��;�5Ä�%׶�8��|4'��_΁$y�ߛ��<n�'�*&>Y����-߯:��*)`$dW:�g|��P��+BeN�� �Z]$j�%ӥE�@Ec! w��]����6����v{n6YׯMQg>s=xFa�T���1N��ϭ	��liWfy�+:{xȢ�g���D�=B��C�=2���n�{X��L;<�ush�k�0Wa�2Fa�/�S.�1���)�kIK~��/��/��	�ç̍�_�nA�m���'P�J�?ĥI��	>�C��S1
��0F7vB��Ev_��K���i�����!�{K+�ސ	�a6_�<#�eT�.���s�R��Q�7���i�Ӹy(f���ˋu����A	��9�"�R�S�Z���,�N#l�I��O���M��R->l��ᅙ���#��{L���上Y�̹Q8FW"���:
���& A>��'�M����M�g�Ƭ����h�f�N�#ü�,��}�]��pF�l1<�%˙�z�\�v�2�� ����b�"��G/Y���#���Z/n\�#	�#�$�e�%��K�a��?O������B*}��W����ӏbf5D`�H�qD˲��6�w������~�q�:���i�H��1�=;���N�4�-M�꟫L����u}��\j�_���t7U�s:[��-�M: &
Yrq����i|ݥa�曃4h�V�w�T�:A��q���/�_xby0+�:f��$w�v���M��RB
-�~o�-&(�K�ؘ��B���H0��q����c��1A���9V�m[׎�.�r����qU��-�eo��UQqk���`�UOOS�ғ@%�g��+���
V,PY~^h#���[�n�f���%@��g�;]p�'vuu3�����*��s��L����k�G�5�)ޘż��M8���'��s���x� �Οھ���.�(7��O�2��377����Ψ�}��?з�;�T�5�*޽�R���0\g�i���SP��ck
���D�]r��<nw�`�ʧ{���E��ӕȔ�4hmP�Er�|�r�(����y��}<��7��rgo;�e�?J���6����)�l�l��&�׀�55�r��OP��A݌ޒ������ ���rEѢLX��T)�m������E=:�������BJ@�yc��p�π�Y�T�D�p��7�a��}|f蕅�N�'԰z�_��o�e-v��s琻�/�Z�g0�`6,H���&yA��qv�}��f}f"!C-Q���/]���\ �ᢥ�/�Z*�t~����] f$���*R��Z�T0�=�C0[�d^\I���1�o�Ps�EQ~�I�Q�kP;�>E��	��)�+Ǯ2,��avr��)�_p�2P_��;�߶65|�G׼'�*?(yfAS�5�$3q�Fk<`̓�����dܝJ�K ��)�6�!�hC+.�{��������5&SW�F�9Ĵ�aO"H�^c7�>��(���y���a ��>6�,�ď��3]C">�$]y��
z�ԁ�#2��j��R�UK�������/a
w�2�/�� �/���/r �F�.}my���K�z��Iں�A3Ok�\>�㎵��<}͎N�dq�����K���d!_Ѥ�}��G���O
��rK�KڞO[�j��dM4|���5����E�����	�_q�{�����7X���gʻ)����U~�1h0�>dZ��m��������9���L�<Z�Qĉo�3'��0��l}���T9aЀ��a$n3\��;<�7hoC�Ve��D3Ju��u�����j-7�?@<������Z�&;���ף��Ov�7#2O�a�9���!�e�~����,�⽨�Wq�[���h6m��=g9rb0o��YxSMT��kw�"�	k��w��@ �G�ɇ a�,�Y�[{��7N �
'�9�O��O�׏��q�©���. �o�.����EKn;�m�":ZTvv��%��C*D�{#W��1���r0�^�5[��9�z1�	S��i&fs|�Gu'�g�\�Ih���X�_X��LG�7ť���ߝ�|����N��<�˼���S-���I�ȯ�\��=�3E�P���	�]�+����,Z�p��NAY��?I�!=+��(c0�d�I�}b<�z���7���28&ȳ5Փ5�󧓁+Kb�jW4��M��4%�Ԟ�	�묟"��I��O��LA_����V���D�@&�oQ�HXU����"�o����P������c���r��q?eK�x�e�t�<������⤹�{�Dg���j����.7[�~�f���ud�>���9����- )��ʦ�G�+��>�9��;�j�E�P۞U�=4��P�d�L*q�:�y�+�8�C���o�ӆM�"B�vqJ�:25�5թ��<H
{�lvӧ�L'���}~"'�r����~	�]B�{ 1j�Ԯ�%5�(���$�[���ڙq��^i{lt���{^ۤ�dcqI�؂��g��5������ >��^��F
�Y��U:-��>�/J����}5wSV��P�� �w��?��k�Im0 A��@c�:�6q�I�t!���~sw��Y�UN�o�h���W���e	-�^p�}��"C�^ ʇ�f+cXA����޻l��Z�Cx�K!9M�.; "o8�t=���З�{zO^R1�I���@%��/�!������Oϧ��2�@�f6}�0��%�f;�Xu�'��G��uJ�� �΋��R_�k��洫c�nE��	��o�('0�&	�t����%�2�el0�ݝ�|7��j"�� ����۠���u8�K�.������sFBы�ɪ+��LF�b��z׼y��`�G���	3��@jtgI��r�gߗ�?=-�õy�oWjI㪜!�N�H��h@��2��Y��MQ�n`b�\���C�PoX�
����0��RHr΁ā��C���� rL�N�%���������]��/��s��E���#�m�����ÿg!%r�8���4��e��2
�0�yr�Z�{�%n�߷*���Y�����?q�՗ӑE>�$����.6�����6�eIin0>�Z2�@�jED�c�r|�-,E��]d��Ay_{)�3Y�2Q�R�s�ZDF���B�31I����Ǘ,ir<9���5x�k�g��ş��==��ߞPj2bm�n�<�:�Z;Q@s�̈́��-��-�r��S�B�1�GB)Z��KY��j����	��y�'�>_�@MA�o�v�$Pn�?������9�'���
��$FR���a :#�K!�I� ���׼�p�+u��	��1���#ԅ��?I��[�E�(�N�7�*��.��N�(A�V-�ui��<�ҏ����Y���͑ce�d��#�F�E���ݹj���'7���q�a��Vm�!��g�LoQW}	��c�(S[�.�� 
��bVMZΤ�H�xg�o�����~�×8�4�r]��FpA��l��^�����ʺ��vN�� ��&Lb�	ȑE�/�� ��!M�u	k\A�����Ǡo�%S�\S
?�jΒ��p�(�}	����A����5�:�H��bDs�����I��o�����t�&~���:>�i�A�&��^����4,����x���w�S>�uxb�A]jKe����UQ^�s�w�h��8i� !�b��l��i�N�a){6��V�F� A����9\q�=�y'�8���|�w4!�\�[M����w%B�|�~�8�-�R�K`RЃ�嘥-��a��X��c>��A��99�M�[���.�2�꧲�lܷ���oDTQ�������`�%qO��z�m�a%���ǆR�G�KVGX��i�#�T?[�Dd��f� ��Wؕ;�5�}��Z3]�-�ۿ�h|��G��SGv<�)�v/�_�8�bV'����O�����5�[��4�.��X<��sS3r.��r�����E�^����t��7��8�]�����u�1"�+�Hg>�����n� �����g�MQF]�&��7Uw짽�b�Gٝ4��a��pE�0M�m�ɀ@��|mP��fI������'8��Ҷ�5fr�#�C�?�Q��ߞ���l-�Z����׻ 5�㝭{��O�R����$ޭ�0rի�c��8�El�X�yjT�ذ���'�X��6�����,�J���y�u���;�_�o��DM���q�1͆��Xh'r�z��e���e��Nf8�É�m�0�5,����%�y\��q�P˓X�fR�e"�OQP(������u����u-�5�N����9p]���@��RH���o��=(�2[����ש��v^,P�xCsњ�Q��Ih�k+f�>�4`���])���	2��̆a������p`#_5i�zo5w��so*��2f\��'3Lw�kw�<��M��a�����K��y)ޯ@!H�CZ+��kҕ=�����ǬWI�9.(���6VH�57���ôۦ8��-����>QϷ�?׵�C]�I������j�/y�#�+Q��/и�L��Ǳ�����*$wU/�R��T���: ��Y�m�c�F4��h��u��N_$��Q��i8�K�*}h4��_�ӌn9D�p��H����u��99����"�F�WO�r�%#J�3|d���\P���@Emq罺�_̻��?>u�R)�w\~����@рU�h+Q~d��?�(��ܩ��?l���m����Z����j'U��ߞ^�4\�T����[�P��9F���6��7þ�����_�uz���i.�>�5-ҫn@�.<26�R{�A���'��!�v�b�2��?a�!���η ����fu,N���2ؗJ���6f�m����	1b�J'�t�M�B�kRH8�D�{��j���[����Ja�j2Y�{�	wN;K-
���9ʖmת����'q��lkQ�	�uo �ͧ��EF����4�:�ֲv��%�N�C˗{R���[۵�OF�j[���9#Μ1/�pS�&������\�aiig<��I��h���MXly G���� S�ٿ��t���N�uw�F5K��;Sh�,4DȪ� ;�3 �[�SZ	G!�+��<����@��IJ�� ?�?�|�!X�j�C7�0�B���C}�"B�u����T��&�I����Z+�؍�R���w���lJ��$�3�fQ��)dքr��<�����_�4&x+'�4F���$J��QAU*���W�o�¢�z��ǭ���Mr���e�_ex�e�t<������$9����R��sju�ޙ���7�� �!�w���d;-����'[n-�kå�<kG4�L�����T�ޅ���� J��;�=�bIP��JL�����5әF�Ñ�r�J,��؁B��qE������Kp�r�<û6�GW�I�T�}yc�!r��5����]�>{����B�#(��L$]ؓW�q�si��!�}��^����0I�e-�k�c�����JnS���@��c���=U5�)����J��#��n�5~T(Sޏ��M��: �����Fk���I��1A6��c�rt6����OK�!�׿R,YwO�Y��T���henW�C^��j�-�����t"�&�^;%n��+�.Lc�aŹ?��?/�1^C3-�!5.~�8;�Z�J��ʨO:��Mi�A�OL�1�z�Ċ�@ x'/π��NF��iاN_��6����eY��1�;����ذ�+Ǭ�Σ�������IoF/��� �	b���yo8�8'�8�	
Ϝ2L���Ͳ�e�(ݘzn6�%H��om�ex ۶0�7��u�s��)�j�w���.��Ѧ��%�똇Ҿ���zr ��q�G7N���n����t�_�M��q7=�W��t��WŤ�WF-�i4͕m�X����디�M���`]9*\&�h˸�^�k����_T���Y�S�nR�6�6�>�צ���;�L���� �Ʒ�U���5�X�'/$�����þނ0m}�%�Ăl��47%��8��\4� �J%j�8z8y���V$?n��*\�Y����LrC���`s�$Z�ˠ�@���'�a��eD����Z�^�[�E�g�c��hm�5�݂���{�=�Y�Q]�Ns���F׹���1D_�cṖ���i�2!�!�x~T�g�4�:;\=8���.W2n�L��;���s��q�f$'�(���b"�S�w�1�Q)��K4��� X�eXS	�m���֚_| 0A»���<�PI�t?:�����4@��p�)
oI=Fm�����u��K\���K�|�I�1�y+0j�	�[�U/�#�ź�z���6������7~�W��¬ɏ�(�uh8u��7k���}���D�%�*��?y#�Xօ� ��ET�$��=�}��&Z�1��X}��Kj�GƘW�:;����C��[ ���YM��C�gviU�*�����¥D&�r�3�oB�])<�p<ʿl�4�ۛڛ��٠�li�ӼB=�>��b0.���/IZ���ɐ\�~���s�����%�W��?M+���i�C�}�}����[�i5z5�H��D���]���?a��ëO�~,�g:�vPi�ZDN_Y������-4�J��Ľ��!t���usF���Ljݹ���U��es�l���d�Ӥv H �n �'Oi��a�/���<V"֫��A�w�ߔ���!0yB�yD��k�wo�p��M��R�:\,B��~��!-�:K;��I�O�3"���q���ǁc�ƟA�Q"9L�[���. q�B��g�·��o��$Q��9�x�G`�/O����[%Ó��᷄��Vb��t��#���[�:I��E��̲h�;Ӈ��-��AL38-N&������BNU�:G1c�)u��� �8�S`'#�O�!��������kX��:.'ێ��HO���3�E>������j����)��e��@���3̌��u�&8�g��akU���}�������~]B�F�2�`wG��	�G �;O�K�ak��m��b�;��|���D#���s` ���Ixr���A^? ���H��
�l�S����F��n	5k���v�O;䢷�@��^L��@�����0�	E��X�;T��Ðp��B.N�;PN�h��gy�Jvɍy,o�5���)���D�w��uQ�l<e�u���'͆	zYi����e#�O�)л��/�0{*`,��\��E�yw�qK6�3Xyf�gy"W|�Q2����H���[�r���Ƈ�~���d]\����R�ꎊ�>=�D[�����r^� y�'�J%��s�[MQ�x�I��k�>��-�?U�)��drZ��a�ؿ���p;��_p�*�H5r��r޿*���fw��+�U3'�k�v�͹������SW�K�J4)�HG!��jC�<�j��0�j{����W �9I���W>�Hn,�7��?�^����5�Qnom>l>���W�C��i�ZF�������#���F�&��m6��}�.��)ٙ�%�wz��/n�Q����� ����
m�2��AⓇ8։�0��i���R�\�D�v���}���ZC����m��ٚ79њ����d�tB҂*��AB-O6_�Q��9|�u`��Tf�1�E_��{_'�U�����m֝�p~��:��{��U��Oh&+d�V�����ߩ��
ˡ؞¹�Z3��eĆ'����Y�B�O#T/�3�6���n2i�	�1��7.\�����zw�u�o!����y85-m�U@�i�<_��a��\.�SB��qv��2D��a�%��V�ܷ�G���	,����-����y�у@m�W��ob�FD��>�MJ1k-�ݣ�.i֗��}�?ua���Y�;E{�ZfNv�
]��9��R�b<�e�q�4���7���)o;�M�BP�EA���#��:�s�v��%�C�q�{�4���.�L���[y��9>�F1��^S�o�&�mY�}L~�,��0Sg���I����N)�XGv�G�GX����գ��2�qr�N�jz��ͬ�1�S����>�ȥ ��{X�3�p��3�	�#+�H��Ii{�����Ds��{��?��^!s����e�0�@��_�}<`�pĚ�I�l�c��&��ՉX�]��+��u��Ψ������A����?4���m�}�ֿA��לM��@�_B�73 r�O�/�6%�%�����U�c�� ohڏ�]0`�2_]�YN��(�A�ôe���x��yta[��Vб�̆u�	�`����=��j�d����7-��(��4��d�����,�bV�-VΨ����G���_ш�o ��17ã�ȳ�Bg=j0�P�F�L�<D��ᰙa�V�9�i�%\���tBQE	q@��ǎ���!�<>��"X�@e��-}t0��~riK1���Q][r{�hG�J�n[2�(��$g~�T�q���iq;�X5^Q���6hI�T��`�HŜ���eg��BK&��ݏq6U0�>��N�J{6w�)U5�Q�S�<S��-��S� ��z����k|�iI�Z+A��c��k6�%����!̛����w
��YVC�e!�h@q�W���8�O-��{�3�s"�*�^V���5+��uc��k�T�^���Ԍ��C��!P�7��n;ֳ��7Q�CKo���=���~O�e�1��X�@�{o/
 D��M��=�z�k����6���������;M��]����0X�+sUh������HT�!�$�*��������{�o���'��	%Ҝ���~�S�e�_Mݓ�3�#���Ym����ۑ��rLXun�ۈ$]!��$D��ǭ��p�ɠ�8�s�ξ�9�z�~���6G�����b�9�5t]���(�-�3�=c@��o�UW  ��-���y��K���t���`M�&�`X y\�.��s{���e� ,T��WS��Z�R~���Ȕ�u��a��VzjLΎ�۳_�8;,�+�S&�/���L5ʾ�m�I틟4 �5"a%��8���48(��8�S�>yh�U�1��nL�m*��Y��[���U�K�H�{��$��Ơ���1�����e?�c�VZ�>�v3�E�8c��כ�(	����z���{���Y(�Q�O�s���F� xX1?pBϾ#�=��i�H1��f/xY]gOd���o=3��T-2��^n�20[;͘Es3�;�#���K�SA̤1 �)PZKP��Z�� �H	�"I��*�_7�Aݒl�l��P$J?up��o�/�ķ�q�
*�yF�\��W�w�l K�dH�:���wx���q+�_�	����#�%�������r�4�r'79P?ˬD+(�����u��2L�J~�P��e͇����#���{�͘��Y�cO��D^�փ��WX���Γ���*O��B=W3�-C�^�Մ$�g �R��DwM����>WUg��y��M���-����MQ���C]�8p7�lB��V#����{*ӗ��y@=b�rܑ��O/j ��T��ɫ]\��ش����}%�N��Ry_?`OȒOD��^�}�%J����@e5P�H�[�D)�óa'��/���}�*~�~gLl:t��iq��-�n� �y4��~���F�\H���7unJr�C5j�˲�gUGQUs�%���8�n i ^��� i͐�aP��3�V]��%��A�����&my]���8Ո�zsw���Ւ6LM�b�`3B;|t~�&�-�EK�o���ξ��������c��A�ò9ǘE[h]r.[��ݡ�b�e�>^�o�rQ�"<��`�%=O �ƭ��,%�Y��<=}���V}�.���#i�[2Q��7#f�����;�C��`�w�I3��a���\�=�ߏ��^G�l)/�{���8�d'^�K���U���B��q�F��.B��Nuh��� 3�|T���]����Sp��� ��.[��l�n��g���!��g�D�&=�����K��������]���-EDw��F��s����\�&���^m!>��6|#�)�YBA�09��。����*r8o}�_?[��gѝ� ��l#����Q�1�v5/ܭqi�OaC��r������&/����`�k�E�$�X��'T:�K�]�k����Cl厢�gJ�^y��+xϱ�����1DC�6�ȉ���7욅��2'(z���8e����W�9��+X0v?/,YQ�E��y���q�e-��Sf��"�ȹQ����@�_�]��2��k�ܘ�o�%/5�o�d]7����R�<�����=��[D��.g����"o��IsG<gQ�p�I^� k��>��o���Z)G�ǿҮ]��aǻ���=:py_�����@5m� ��i�*p��f�]���3�<k�R�T\����vܮLKQ̲)�!>��C�,R��˺V�Fj W�H9dP���eHICF79�����`���&*�>��f�5�%�`CӤ����˸�R����#cͽa%�%+`�;��i�����	� 
,w��6/)�P	�ۤ�0 �.E��mJ�Z�<�ꇓc�������N��������b}��3�U܄�$��|��ٵr2�#��1�Ưk����<�Ol}��Z�_(|Z_	��m,�l/�E����6"_��ⲵ��+��m�ʻ����/UO��h!%dk�MӞ������|�2��YZΦp�`�j'aE��+�j
!T�`�����2��,��7y���uƕI�u���]ӳ˴�h-[�@��u<��%��f��w뱁�)�w��vS�2�fEa�K���hJ���љ'��,�.�dH���]��l��m�H,x
/bab垪шM��k��������S����a�F�Y}�{z�N�C�
��9��t�`Ȏ� .�q�abdj���ov�U��ΑE<�~7@:C0v�[�%}ݩC�8o{ȩ�ݑ��i��oê[4:�9Y,y1%�S��t&�����̙�]g�t:I���ɖ.X"��G4 �V�y�V꿍ܮ-w_N�E�<��v��Sށ��bi�Ƞ���֕3vY��3�	=S+��-��7��AK��?����G?LD�!�y�9�&0�^��8e}���kؐ���%�Ϭ&�=����8�+��Ǎ;:7����E \���Z�l�\�E��~��02�rso���B_��)�4��j~A��TF ����U`[S�!�o����I�M�z��Ⱦ��!"ɍe��x�Ũt��������Z�������x��j�������7l�%���O]�d1��z9�ϝq-�Pf���jG�=��֊x=���ѣ֓��Ohz=AP��9L;�m�k��|�/m� Ҍ���B�vq;d/C���Iْ�<�g<�~2��xy�{���|�}ogu�r$-���]���{�4n��$o�`�(��N$¿����q��i���3�N^�;�5�I����!\��&�1	xI8N��da�}�*v�U+���O�|J6���5toBS�	�Õ����� �@��Pz�k7�)I��A,q�cnB�6"�����!�;��Dw�!Y.���/h�!WO 9����-���ώ��"PN"^q;cd��+�/c	T_����ϧ���C�j�!kkit2�;�,q��k��f��~KN��f�O��13=�Ā�2@���/E�`��3������`X�q�96�5a�[�lr��;W��������Ue��7#1�����~]���ek<�?����k�o��'a��	@F}�(�YUC�e='*ݎh�$&Pқ�)3�_�[�5�l�z�u	��㳄-j'����x���C�N];�|z�5��~�G�)�:F��T��t��s����H�=�Hϵj��W{�Ī�31��N�c��oEU�
M8M"��`S�\��w�.�[��jX�{�é���Q�R��
z��fA����q.6L��ȶ��V:��0��N�/ڸ��Ծ�gms�@�z��p/�%C��8���4�oC��j��nn�y�՛�n��*���Y����7��q鑖=�$P���qFD�l��ve:��A�6ZI�░�*E�bc��-��V�k޽ӴNRr{ZŏYCQS��swt	FM��1:�A���SEi�~i�`nx4�1g�UG�p��=.Zl߯Kq2��on@`�KM;�l�sT[�՜qM������S�@u1 �)���K�Ι��ڛ{�	��j�8�S_��A������}P�1/?�z��Q|�*`}�&�
�>�F�>��&�AsK����J�r~b��o�+�u�	��K�#e�a��Zk�,���jn_g�7���5�����(���$eu:l��-M;����>|�8'��X����#X[��r��ν{����X�"���ҩ���W�Ε��r�=��W���R�y^���6� �-���hM+�9�Mg,�~��%�ԑ��:Ֆ�((��冚]_ep2�l��S�j���W�b���r&�����bf�J��̊/�n�jk��WR\�Yr؏���Qh/%$��M<�?�q��
�(�y6}z�ݛci%�{�5��$H��D�@߳�Y���?����#�~�*�:��i��0��)��{�4w�Q�z����1*�$�uinvR�j|�O�&MBU��ps���-�	|� �s�ϋ�b�i�a�a��΃��'V����jaA��s�J�v�KK�yx`�ox҈m�w���-��M��C���:B�+`~��\-��K�׃���i{����Z�iF�co�A�U�9Bn�[C�.�3��x�]ŷ���ouEQݟ�n��`hU�O;�>�%�?�Ǘ��x>gV�0FjL�#D��[m�o�� ��D��h�R;I�
���S3�?�?��9V��8&����G��)J�]�v�8k��'�K��Wj��7�F�����.]�������3#�>�C����Ȥol�+�&/��K��Cީp���|���gO�Z�D�����-�v���8�]xi�(��w�=�ʓ�*��1���|��Um����1~J|~g��`��K��i1��[
��^�r�Y���?����"z��;j�l����1��lkX5���lrO�k�-�������=��l�b㦤�E=�~X͕0T�r:��m�x:��1����ݡ�J� hy�M%�z�lH
���D�BB������z�҂���6"'���z����o�etW�ߢϻtX��C0qtz,�%�� �y�0pq����K>f��"�5nQ��᧾GO�M��]Ę�=G�`��
�]�
�Q��Ry����$�=��[Z$�J	��V޾�o�]s=�Q�I��!k���>1�%�u��)��d�S�(a⾣���p�I�_�j�KYF5h�K�(A*+�8f�KH!�63ݹ�k(O��������	�Kn�)/�,!��C���gY��f���ԟ�k�Wz9�9C�M�zH$z�7tǛ��a���S��>�|���h�+C�奐�����@/#�|����6z�p��^�_2�-Zw0|)/�[�$�x��^ _f
;�m�G��7���Kڦ7��O��HL����"���}9�ŐP�W�bA�7�R���3ѐ���d�]���`u8�7*,O�;V��Хt|�h�����秃�E>�����_��/�p��\2���b���K��U��h?fd�E%�Y��-�������W}�8n�ZiX��[n�'f�������T%K����g�M9G���'<�7�l��Bxư;qu��}�8�����-��L@�?�<a}������i��4ݣRq�v���2zY�a����n�Q�`�B_�,}P,�?�����B�+m�Y��:nb�
�ńUM@&�k�٣�/Gdڦ�/WlL4���a��Y���{U\UN���
��9�+�׻N���q'/�通Oo�K1�xm�E7v����:�'v���%���C�C{l��,���p�ʟ|[��9t�31�S�S`sC&R��[�Ԣ�r�gmg�I� ��D$!X��<Goػ����)��,��N����^�Q��Se`����ț<��1��31b��S�	�+o+sN���%m�� 	�:%�1x\?�%!��Z��"�0h�{52�}r$��f���D~���&4̐�[��w+7�͍�����������{�T�u�u���j��D�5@��j�����_����i���J��,���L%��U����
�mo#��ӏ7�h� �Oc��x]�ze�eRx�%tt����E�����d�۰�<��ϧjF阙��7�!��R���j�d�@��Uy��ج�-�������GEAƚ�rc֥�ȅ'̣�~�ۊ�=�+�P���L���&����i��/�|��g��9lB��q6�c��k�P�W��<4�r�ع����%`�}j�t7yr�.u��-]�<{� e���C��.(���$!��M�q4�"igJ��Cu^ǭ�Љ?I���|Y��Դ�L��*��c���{w�Ś�U&M>����J�[��7��5�QSo���j퉉' �����\�k��-I�wA���cI�J6],{� ��!H��c�Jw���YI���[��h���W��T�n;v-�x���"�^����5+Z�ycD��ŊQ@�ʋ�B(Cd9�!���_;����:�y���y���R��OJ�<1N�U����@��o/�^Q���w�0%�,i�6�A���\M��;��s���e�����ޠ��:h�>ɦל��@��wA��{UoI��'ɝ	[�М���4d�~�Ve��݉C�`��Vy>N��ֹ��G�c�u�̈�"���j�_ɩ���lɖ;�)��N�zC�c�yd�GH�=���+�o�!tSc0���3߃�=�q�e��W�v���Z)��K�ޮ��J6��EYM�-�`N��\7���J ��S���$8Äo��iYR��}�LOx����T��jL]ȑ!b��\�b���I@�/5��¤�/`Om�n �U��ë\�%ޝ�8�b?4��"�{�b��Dy^��皫n� �*-<kY�ʷ�]�:��NΑ��$�1!�L�>��`��2!+e5���swZ�:���E�wch~�������}�Z{��Y^�Q��BsRF�e��9Q15x]�t*���ҕi�����y�x��gŹ���?=)�m�
��2N�Dn1��&��;�`�s��1�7����R�s��S��)1;8�)F��K�m\V/��6=�	����3�_���A���b̳P�{$?�����B% ҷ�Џ
��^F�@3�Ma��6Ke�p�}�m		�BZ!+a�1	 ��ƀC#@E-�+����� ���|�7�mmPϔ�:�(�,s˽u�� �(nV� ߝ���.S���}=��Иr#� ��J{�ɩ���ҋ����M���0�	R:�`�{�8��W�R�����p��d �y��N�.M�Ȏ�4;�g�Mc�[���ڥ����� Y�]�(
p-Q$l������=�ǃ�� 7�MȐ���~b\Q���a/ /(��lh���\���j�ǌP%�I�H�?��?�Δ[�}��=�>a�Ӷ�5K�H��PD߭Z��r���o͉uɵ���~�(�:�gi�e�_�V��-j�6�)4�e1�UGU��:���@�ud�����j7	��AS�U=ĸs��Z�TA��� ���G�X(iS�a��{[UV���[q�A��Zߥ9���y�<��;�H��w 
R���M����K�AB��O~��F-�<�K�yO��y�X��at�ĵ�c*w�A�9�c�[��.�ss��X<��rqo0+�Q�<����`C�IOvVc���W%�E���3�8V��E���#��[�ݰ�m>F�����<;�%'�mei3ɾנ����g�3�H�K��Gb�{)e/h��$C8F�'Է`��]��ug����򼻠.xV��D.�y��3^K���b ������1�R�AH0�$�s|�b��򊚝r����g�]��l�ګ$�0�QSl�9��]9��#��wXP�N�%EԵ��9��x��mW]�,@|�Y9�ϝI�f���!�6�Զ�@rnd7��?���B-�VJOl��c��ק�5<���g��O����?��`L�l��G����]�E�ŇXȉUT������������\7�����fJGL�y�ݷ�H=�'� �ۢ�D9��~үJ�m9����m'ނ�z��d����e������7��2fa4�0l�A,r��d�yȧpq|�����8f>�,"(ºQ�������yR5�hMYaX���O���&奎�]����	lR4H�q=�5[5$v��u��@�hL6��s�]�Q�<IT;k�Qp>l�O�^8)�()�u��ӻa����*�p̟_!��摆5c(�׃�q*���f�Y����3���kck�͊�?����dڛK�/�)J�!4��CrIQ��O��6�����W5��9��*��_H��87��7�/��ǚ�b�c���>�K6�+��C�CI�A�+����"C����#�rV�y���Uu2��(V��g�pDw�\/�I?)ݤZW :�9E�Vm���2�,�I�;�a�������:�Ճ 7Xk}�
P�Kn&��Z���;��H=�� �?m��%Ղ�p�2�UO"@������|P���|������Eٟ���$_85=�+�̝cnG�p��,�U�hyd!����Y�H��}n�2ɷ�s��Z*<�Vs�'���ߊ
��8�T�U���,忈�o:K�"�7/<�����M�u�����*�k->�\@���<p[�>ҥ�����\�-!qv�Oj2l�a����g�F�ZS�]G8,�;��ԗ6�U����m��b.�-b�����W*M�\Zk��/�0�]��+#���p�]a��Y`�{0UN'��
.d:9��k��s���,q"�DXݳ�u�&o�"��,�E2��4�	:�	v�c�%s�Cq&{>N&���i�w�%�N[�)9�
v1�qS;%"&��;�N����G��F�g(z4I�j=ܿѿX�,�G�л������Ca����N"
4�2W�,�nSTh����Ȗ�EČp�3�o��	3ow+N���3��w��5�1�� �?O!į��/��0C��pK�}eJ�a`їZw�,/&O���4m���+rׇ�qq����_���K6������R#�i9��po��������_S�d����6�����2�=+mU�>��k^oyw�o)���N��˹��3|eRR|x���tryGㇰ�m�zj�ۋe����j�@G��e7"�*���х�d'���0�>��-'�i����G�����f���<�����������=;YP��L��A��b���@��ܘ��.�t��B"��q1�����ǿ�E�rj|<��޸����yV�c�}e5�ύr�P���^]�p{g,,���,�(���$x�ՓC�nqO��i�����^@�kc�I�ٰ�׷U�yG�gG�?=��>����`߱U!%(�u�J�J�R�5j
SJ8�9�r�$9E �f��_�k�HvI�	�A"�$c$�26��Y���!���!�w;�Yd��֛Mh�9�W�|�	��-�;��Ddq"��r^���Z�+5�Sc��%B��ŏRԝ��C(�!��Dj%;g~�6T���^�t�#���&Os51i]�vu�@lG(/�=���g��������m�6N��Q�(�e;ͫU�.ф����< k�0��U���3|�V|��5ܢuZ��o��@'��	v
̜b"�e��es݄>�ںj��i$r�Q���"��#mu?~��Om��T������e��d���z��ʩt�	G�O����V���t����V߾6�=4�O�`Z�W1R&�C�����p�Y�s�%Go뀅�MX�\`I�\��ˤi��\�qQ�_+ �?��RO�E� >����ג8幧�L�ԙ�l�˷̞!�#ߍD��/�Q7�}���J?�mi1��0
���W%y��8��m4I^"�60S���Byِٛ�W�n�X*ț�Y����{�|L��̇Z$F���'����Ì���e0���PZ�x��ǳ�E�5ycC�)�T���)��f�cp{��aYy%QI�s-вF���I�10,���]ćnq�i�JR��px�7~g >*Ŧ��=$8��e�2	��nL��4;^tfs�Yo��>��"1�·LSr��1V��)�h�K�,������	�#���_h?�A.�����uP��)?&�K���I  ÷ܯ�
[�F�b���Ɔ�K�KHM�ji�h�k��d�+�	;��A1�#I�f�>�b�6q�!7jN�k�U����(��RT��upgf�#�m�[?��3n�W���6뫮�#����LCv�ĵ�t���Ș�'�;�Ȭ����V�D.
��G�3bWDT�t6j�*���U c��Ma�e�/�Rg�.(��
�\�0���5��[K$]�b'p(��lS��ۇyѹV��Xs�(�w�*�=b� ���/{f煏���+5\}���Eg���X/%Z��C"b?q ����ί��}p�i�y/���X5�_�H�e�D:;6�I������4��f1~G3:EM�i���������U�Qэ4m�0���d0�Z��u_���j�Wv�\y8U��,s\L��u?Ӑ D�)���aid*a�A��VSV���A��� ;ۗ��|y�8�eW�#g3w[T��c��M�Q%�-IBl�C~|�-�K��׃5b�T
���)�E_c��,A+�T98y*[�K�.�1�xcS���O-4o�0�Q���dEH`HO��/�t��%�k �M���?nV�`-`��#��[�Sf�|�����;�6i@��[�3��p"V�o��.~'���G>�)����lf�8!Wi'Dy��q+���ӟ�D��w�J.���ݿ�|�T��3�⏕y�����%oq�\��\��韁Waq��r�8\���,gTW�����|R�,�U�ts�]������w���	�w`0`�'EKӷ�=W�*m���'��|4l!��3Ɂ=�_��z�5�Hr	�X��xO?lD���+�qJ�l���>����w5׏��b�
Orᢣ���4K���ի"��7(EsƨXÝ�TKya�|�u��ƴ�'����f �SJ�J�"y�^����;���c�D��=�Y��X9(���j'9l<zE����ue�������,��u�0g>�,j.$�v�y�>�q�t[���Cfy��"�n�Q�Or�Q�E�4}?��Ϩ�ȗ�|����m�@��]���t9R��<����=��4[DW��z���7>�#�sx�Q KIϖ�kru>�����K�)����г���}a%��сp��_\������5^�����B*�Pqf㇒��3��ck���%G���4�ܿ�cK��)e�2!���CM����Ҝ�*��l�WΎW��9��z�C��H�G�7�Kȕ�t[�g��[�A>�:j���C�\��Ƙw���?��-.#����S���#�0B$�����ת���w���/ZW�Z�	��� 6��mݡ�-���ˌ�I�Տ[�>��㰦�r֝}oPҐFg�5s�����Nц�e�;��`�S�����-��O}���L����|���Wx���sEt�n����_��
��4�����x�K
�g�}U �h�"d|Xt��p�c6��~\���➮�
Z�V�Q��'N[�Ek���fT�Т�r�Ã�էƕ��7�+�������u������d�ey;-�Q$@敃<�u��7����1�~����4v�2���a}}����Է�J��xOm,sG��Xl�q���=:�m�����lb�u��JM6��k���k��˜�G"ck�+мa5��Y�+{�Nb�u
��!9��A�q��Q�q=����ʀP'o'eͮ
�E-�珫>:t&�v%�#�CLM�{yP_�b���쀸 [e�9��@1�8�S�&����^��D��(�;g��I
�V�:�
X��UG���'�v�/�����^P�N=W��o,DS�� �3��ȑ�����3��n'��	��k+)�_�5b/���0WQ���?}_�!��"��_W0x:��n}����\����O��&j��u.w�ɨ�+���=3���o�V�c�n���_��g�D@֫��C���|��_�c@3���B�"���*0�x�U1��� @�o���Io��{�E�x˔�!Ә�e�^>x�E�t���B;��8O����<�f:H�)�$j|�����I7}��ȿ�Ѡd�d�.�Y��N�u-���
�G���K����@��e��g��� �l=֦yP���LL�뻜�P�͏��%�����V��n
B�gOq,h!T��z����B<*w���P�,I[��}`��*trU�ɮ  �]�8{BXó6�hǬ�(�N$�C����qjR�i]�ً�В^=��]�I���2�R�4d݁���oK���֦��CU��`l�Jg.�mQ�5�tS%0��t��� �)Q�a�mkh�I/�A�j�c�ij6Ӳ��V0!�CE�oww���Y��Q��h���W [赤f}-��dϟ�p"�ya^�̇�mf+Խc�����R�������N�C�6�!����� ;BW�qH�ʯyt�o��r�O��1�P���i,@G˰/�<��U� ��k���^���6
;��V��5;�+��"��u��DT��p���4���0�Kʢ�
���Io�$'��	��o��78�M6��e>�Ys55X���3�����ڀ���%^9u��5��>���J6�-Q�Ɍ���ߍ!��R(zy�)�o�HG���ky�R.tI����z��w�=�"��[�rW�MG����*��ԑh� x���M�`D\\���_�����L�:Z�z�oR�	f��O��M�Y��

Ll �G%���͵�?ک/��^�8��e>�m���<��!�%��8��84�B���g����yT�]��4�n8�J*c�Y���N �7jd��\k$���~#�Gx�h�
e+��RNZz!��sE��fc�ϛ���<��o�c�Z{� �Y��:Q���s��F�w���1+ ��*���)0#i���4x���g;�)�A��=�$��f92�G;ngc���;9�s	��m���k�)1�S-_?1q�)<X�K{�̃��l �	�6��I�i_#��AI/��X!�P�o??aj�"b� P�7��
��F��_�CL9\��K�嶭�A�c�����+�v�	V����#�����&��C��z̼p�7%O����0ٯ(c"��w�u�������o���и�s���>#	�U��[���ቔ�<���I�B|�C^9�x���*����J�.Y�W�*x/ط�ʉ,�̒ >q��ġ6M����*�_g=0ͺ�@H�%~G��Kùl/��]W]0��p#K)l��I�B1i�7��t�ln�e�b7�&��t�/ֽ��@����"\��P� �Y��}%�L��>E�?̘��;�E��E�}�b���,�,)�5��H�SpD��q���40��k����I�~S�:�Ri���Y��Z�šl,�4���C��H����uZ�+c�j����w��U3��s7I����ڮc ���x���_i9��a��1!VIr���Az�<�[�]�|yJy�T��R����w�����<�M~6���PB'�;~,��-���K��o�pף�:q��~�{�z��c���AF̅9��y[�0).GT$�I �NK��7o�VRQ.�����`���O�LP���%���Ǩ� ��V�(��N�#���[ꏽ�����y�;zr�[mQcr�3jaM�c�
P��)Z"�K�G�)�K����s8���'J�E�(���ݣ|�Wˊ�2?�.�H��:g��/�3ԙ���C������ �\9��wk�y2Hp�ZWN��e�)g`��*J����WO��@]I����w����~�{z����ӒҬ�~�m��*�"�_|��I�EybɜM;��Z���aD�p��r��Q��r?ǡ>�S4Mٌjml������ֵ5rE��]M}Oͤ��^G��OVʍ)������W0"E��X���T�,e�7��ɼr�����O��NsJ}C�y�A6�ϝ噱EPD/�-�4㯓H+�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��} ��UWP�Hh1�;�f��l݇�Jߚl�.�u?W�������Jd�WT�VEk_+�o�y�wϢ�w�Yc$�����^�l]b���
_��Dd�3ٱ���k	�9%]���^Al����}���V<�
=��s�'KK9�#�~v����B�I<���[�z��!������c��D�P �=�����:����e��$^�]�]��.�(� ݿ�E�o�hO��z�Sp[�(�혾��K�Ǿ)J;ǜ�zH��z: >ߌd����+|�"�<�H��l�
�M�tc��X,�D��e�b)��n+yL(�f7X2E�3�.�/���1��7��؈MsQ������{�+'|�.��C��@�7_����i�)j��{�!� ۷͖ٳ���U�!�0��\���� rbExy��⵭��T�cUc� �'�a6&~lx/~"\�&���+.G�����k/�~��<�Q�]���/�UZ4Dn��&]�\ֲ	0���+e<�6�p����ꓭh����@��#c	��N�
N�p��Z�(��xmW�wyM��({Cn$�]x�I���b
�^_�Izmh� 5X��.��,���$J�K6��\����ᡊ�J,+%��� ��^�����Brn����WwJaÍ���>\�D����Kq�Ţ���c���"��Y�P(�=�q�#�2n��M�I��6
���d��!N_W�q\[���#AC �+�IR��<R==�b��u@������8���,�B�u@���zY��Faoo%�/�0To7���t�.�Scѥ�3��[�>f\�x6�1�KK ��z?��Lh���	��[��� ��x*l�M�5�2UvF�h.G����-�+�Yʸ�w2��R޶5����tze4�l��(i4���·�2'����s��sT�(�=Ĉe,
��a��]���|���n=����R	���v0��l�i� �.A����:�q���ǅ��Gv�3V[�
�H�|�������q�#�s�H�[�4 ��\��d��(`��]�:�ŎbՎ-��=U*!�c�?��D_b�=@o|np�Fw�.���b�*C3����8<y4��Z������w�l�|�e��B�Y�Q��'d(��rU)�/��TH�����vٶ?5e�Q����>[#�=��<�&+r�R�>P����Ṁ��/�+��T�������ǽ�^�y*�1XX䡞j=bU����yx��f�ҿE�0.�����M(q���s��&�*o{��*|�@�.��Xo�k@�y�_���b!2)��~{tt `f�B���DU��=�\��<�����y7���aG�À�TU� kM'_��&��T/*MɰRO�����G&��J��q<8�]"��/�l�4pZ�������}�	�T:�?M�<Rlb�S�Δ�x��t�e-q��6�	s��Nט���Z�%�$\��=�9i{o�&�����u͘�i����L���Tzh�P�5��-��U��}�������a����w����& J�&�+Q\H��]��lc�6$��n�{���_�J�i��O�\Km�����t���p:����֖,���()m�q�8R2������I1m86�9�D	��_�Tq\g�:KC��x�K.�6L�	�<�D�ߠ�8�./��X�{���K�F��Ӏe����\C��%�Y�f�XW��}E���P�I�"�������s�%�\�U5�},������<�逿�+�����4�Ā��c��'b0-�E�i��b(Q����9��٦�3�dǲ+7�5��GWx}��f���{4�4�� ����*��P��s>��Ef�l�K�_x%~��:g��$ a�-�H��8b�q�i�����Γt��&~���[R�ƕ�Jn��](�Av<����R���_5�D^G�Ogn�����Tzu�,&K��Q��t�4C�w*�g��"l�]y��Bk��nIA4lM�Ot����j�I�{�σn�$/��A��-����G;����0��8Γv��1��21�DW�( fN��#߿�`�m�1�,D@:�oX6��n(f�oM.�^�S��1����Jcb�����]��\=��[�&���P��n��t炱�;I3���Ռ��s����ԩ(�!@d�`����1��jIߕ܏?}���n���Mn2�6s����5�h���{�`���T)��*��t6�e1�VHP��g�~���|�1�v4�[���Ϳ����C�]��)��;o�0��ʏ�"}����s$�
���]e�5"��/�J.�7![
�*^�MO�����ο�F{/DU
�e౞7e�<�b��3��
����c-D�Y����^֛��|���N�b���49V�)X�I�#b�]	�A��{���!�!X��g"ϩ-��	a�����=p�;�=�ה�����)0��=�4�!�L�֔�Mm�RF=)3�BY�r��΃H��#��wy���~ �	ZR�Ʒ㛖d�>0�魬DMAͼRs�o!	�f�%�_�0�&Cy|(~:�K�Ω�Q�@>�{������g��yy�rվ�|K	E�ʘ�S�3rTz��T�M�;(�7\`ƪ�u`S.�G��=��N�d���-u��n��<`�w�S͋���Q�6��I-2�c3�-����Q��r�]�8z��篈�6����<�q��hk������5	UI_!m�EYjy��{E��ˢ��3�޹��������0nU~&������&�mҳ8O�2�
&�����P�vn�8}S���X�w�Ρ���hiy�p��`�@�Փ^��̅���z��֯6��Ã��?Y�Z��۹*o�"�zjD/ݎ3Z�ǝgZ�f�.o�����C�"]+����4���}́|s����n�o���t�����{ ̺kI�:�
S��|�i1!� W�6��G�ր�,7~#�I^
��*���>z�A�7#��$�Ϗ֔9��2�T���	��0e����#�L���A~uY�4�$����>�c03U/U�X�#!A����Xk��y�: ���ϱ>3�Q���9X�ϓ�(79�<yX�6�-;p�\����)*�Kߚ��%�)a�h�P��i7r-�,�������v��0U3�>�����4�s����`��8>ŋ9�;�M��>��##XTPゥo��˘\P9Ҹ*�2J���N�����1�eՐ��dx����hk.*����Ǯw��C�T��ek&*)�7yr76��?}���z|�cP7W���ҎpLb�Xm��r?ua�D ������||NR2��wقL�	��1ޒ�1�T~ަ'o����G�^��fN�j���2��s�u�[���Pi:��g� ć��&ݙ�� x�xE�����*"'g� bȷ%�1��������Z��1;��t�E5�Uϟ���*f���Q�(��Z���Url<���`��I՚s�����6���8}>��_4^B2-��:�Y�{FR�%i���o� A����SV��҆M;[�${\
�o-�S8� .i!?Xc�h��&	��[e�������$l�]5�<]v�7h!�ߍQK����<Y$,N����%-5���\�HX�#���W�����*+�'��Ԧ� s�-�K=��
���aH��k�����\h.�&�q����W�!��v�V�?,"�S+�.���s�:Ӿ��u��vB�4[��Ɉ{"ɧRFc��6�qp��&�JH���s|�＀�%�n޻G�P�R�mX�b�����]*�W�6�E��%b'��ooN�n��wl/���y;*�,֏~ �<�V�ۙ �:եلw�pK|�߱Ɏ��Τ�Q�d��ZI��0�)F��g[:������XE?��Q)�>�Vm#�>`����+�{p,�P�ޅؽ�DFq�85`���8��H��o+Xn~�`�D}҈�<�w�ˎ)F�c8��]���ʡ>A)A�ޒ���s���T%�aE�����7���mx�`�:�������!�*C����(`���z����$�1r�p���'�=z� �I�>���~8
e]�%|F�ק@���n���H���Į�
�[2�x�S�m��F9�w+eNeXfA�w�B���1Aؐq��"�/߫�m��-!m���Ơ�o����[2+�������$Q�ۦ��m��'2�?��S>�DG�ҫȪ�.�x+_�ؒ���x��;7,��#��+n(���_!l$�)���.:���/w7�ܸL�{:�7$��EL�������i����f���vmǲ7y�$G��.]��c)ŕ@*�~����@7�ufC67���y��B��[L�̷4w~�B�c���%C��=|�.*�y�� ˔�EP1q���� I\�W���.�5�$4���j~��ɱX�2&��ϖԥ��j">�w�(�v���� �42�e�}D�W��*����(�hoC��܄��o�6;*wv�Y�k�;B�^�13�O�G��,���G9!BY{�����+y��s�3��4^�a�=4�����_'��@����6�3������� �D��4-֥N��h@�e����v1(�˚i�{�t��?ҌO0߂g �D,��۾h{����!�7J��,TKo�O��'�v%����п�9J��x��a�!�o�<dl��b$�����גe-�cN7���v�����]���$�a�u�����t��N!#3N�_`p�"���m�I�'��{C �Q��ݯ۬��ur�����J�3}�ͫ��:����!�iV��+u���:g�_G��FYdO�ֺ�I��
g@�`�j>�1��\�@�}��O:g\T����B���p�)�?��>\ݨ<�!��gy���zٶ���z��)��n�%�����z-́���Ͷt����	�=��\�u5���T�	c|�,!Um�����'���㹩5HS٢���e|j@��K0T�R �����A�Ϯ�A>�Σ�8�zyj�B�ϸ�T|.��d�e�"��]���3C����	��HH/O��>Rm{�D�i�i�VI�5�)�\�{�S��+C�֠,c�r�i�Dk�ʱl��8y�?�v0{�OG,xl��Hk��D�
�ؽ�״|¤�EMcP��)ex�5�T��
D
�i+'>��2ٳ0�E`�0
l�=I$�ҁ|P��6�G�#'d7�h��#�ԃ��,��M:B�� �$Dq�q$�	����i›���,��Ѥ�;�pF�XX������z%���>�l��e�J�����W޽�k �kߊA�(9��������r ��ۅ�XY�D%����J`�⏈�����+�R�rM���a�:�cm�;"��&�r�_2�xD~6eI�A2LU��:9a����L��]�c��q�Q��ח�v?��J�~��YNOa�?"����c{9�D�&\4G�*�b�UO��a&�O���E31��2&�;��<.�^�Ec��C� F�l��H+�t�v;m?���k5�LC�+��xV�ߙH�Pm��#���a9k�J�V���=��0v��bm�
���3Wp�F�j2m�^�S���@[�C ￟����A;��	���t���!���;�}���-Xm���V�N �;}2�˛�HrY���M����hS�t��V"�;p�h����k���RQ�9��n�-(F��fh-��IP}]�/��,� �����B�ɼ���
.~�Ѡ�}(2tB;��O��NO��Wt���[
6e�o�h������W�d�o�o�8Wy�{\�M��(<�)71������dBH�	��u�.���s ��)UrDW�1ᶛv
�
�/���g`Z+ʮ�����`����y�P-�i����{��&����]��_����B�{&������=�۪	7	��r��S�����������vͶ$��@P~�rq��ע
ڄY��#���/�^�L@��Du��5�P�r|�?��ZU��nq��^@��=��J&5Ir���Ùf�h�<�|k4s��'�;s`��tQ"�&����g8>R$Wkn$�b�!$�s��h��tŭ�̠̄�M��뎄Pp�/إ�";Y��Fq�T��D��3�M3#��N���(գ'g���.
����?���~%6�©p4O\Uo�'<ɾ,�M�y�,`����Ms$��9�4��M�
���K>�`�}����}�\�#F�1��#�}R��ɳ9��x��=�s�ZU��ƿ�
��Ή�����`q�-���섥��]|���d���z��5fz����BxR#c�	��Auz����`���I�����}�B8 �C �T/B�����̐��Ų�E�6��4��y +$/i���*�%,�X\�AoD`.��.���y�W�	�i�����5�;��P?�C�O�D��5���L i�'��GP0��V
CԐ��_���:�T�eo�A2^�ЂPcu�#��wAؒ���s�y����Ė[５���!���x;���^7<��BT[�YR޶s%�����V|����I&���ѷ����@cߩC(ĖWup^��G��Oі�\tQ�R�]"E���g�dQ^k�C�*Cp&�n�Z�����Y����0��ߐ��E��8���+4���0��w�J�z���/����J����J��bWD �V5��_��ij�.jw�c�$��z�٤PlMf;�݌�_���d���N��[�9�t���l��-����������߁'�4�9�K�~f$���Ċ9����_K]Y��}������S.��4�, ����88��j��|�e{4$N���M�w.�.y ̓�EtZ�X�DՎTz���[��V툶^���-�;���|:ǌ%`H4mz*,?�|�t�+lg��,{���=��j��=�SvX����=WbWG�^�]y<:f'�YEz�.��j��Ρ�����N4sAN����{�k�|�B�.��3(�@�T�_�&����)Z�{�Q ��e͆���JwU��6� a�L�O���GRe
y���⥉?�D9U���Ķ'��<&n>I/n2G��5��G�4���� �nA�<|�]桎/�U�44lQ�E�L^	 @����<�8��`����� �X
���{���M�	�|6N�p��`��Z��]�hM��gW��}��{3�e�����9)��v�N�{�9Jhy�5�!��8Խ�t1��jh�;:������ܢ�HtJ	��+�K��X��N�ڏz ��2�З����>JQ/*�}vh\�l=���`�;UQŒY��;�����I��(��q�;@2^P�=�}I��06�>�����m�_G�:qLc���){C����^��Kr�L�;���&��S�|�/d�vX%��K+T4З6���/d\`%.i6f��X�ݴ}	�H��,I�\=����U.�%!p�Hс�� ��f<������M�uM�s���Icû�kZ�-����q��Q�X���J�����(KfU'[��n���t�}eڐfPM��?T��QS��ͫ�6*K�~��-�D��f��%K�*�xi�'�����)�a��)���8&^�II��FU�G��W�e�j�A�ŰjR��� ��I.���"R�Yw_y�(^Z�g��6��T8h->��,jz����t
E��;C�g�!&l��� ���}IpAx�Oc�Kt���n��.�ag�K�)/�`iA�������__y���:U[��״γԬ���m���(d�2��+�^�$�m�^,���H�Y6Jԗ(�ԽM��p���O���ӗwc&�r�K���	~Ǡa�j'�S��P��M�Ө0�F >�O�3�H�� �7�?�P�a�m��!��`n�%�uG�j���k��RC�n��uM2(�6�TA��Ht���(�D";{>�e�s���.b���6+6�z�H���g�:;�+�x1�3��������Od$���&]�>՞�{��Yh`���e"��K���đ˶��]�NV"؀/8��.��<7e����!����}O�1�.�
ôD�J#e���7J�_<��P�w�4��(?�h��'�OD;�w��c��=��@�_���/�ȫ/�PVGy\�ȱb��`���L��f��b��3���Ҿ�m�bUř�^x�P��pqQ�=����98�#���x��m�ZGh��R��3�]hŶ����_��?x{��T`��A �'kRZ����:fd����Iଈ��̀�����~�*NJ��9Z0�Iy���:�x��NQk%>1����fޑg�*�y�񆾹�]KM���\#�S1��T>��"7�exz��7���`
/9MSrknؿ64�5�dQ�-�\�n�P�`ಅ>�c'�QH�Ϻ���'f-4��E���#��n��t ��l7�E{P AX�_�&k�Gm�e�5�����1_sY�k��ߵ�������pZC�����c��8Nn�t�ϩdb��p�&�� �|�2y��� [���n�2�Sv褀������!~�i=�$���@~\����I�ѕ�)��s������Z�Hk��8J"}gz_�!2zZWӸg�d�f��;o9���I�"�1���A45B@�A]�|�+`���mo�gYt��~��� �.I���
��|�!D�$�5�=h��F7B�I����JI�8���#�$[����K
��#L�)ɖ���0�Btѱ�#Ϩ���u��a4��3��>��0w��U`����K�!�����qkX9��~ۨ�a��������
��XH5��lU�� `�z��;4*��������׏��܍�)�'�h����,�r�(��8�t�X�v�SgUڠ�>`⑟J�ֱ�k���?9�+\'���}�u��1>\"�#��JP'Njow�)���<9���v�Kci��[��(Pe`+�(���V<ý,$#* �M���}�7��D-eL>*�d!7�&6��?LR������W���0�"��N�L�G�mR��?�:�D��Ƒ��j�@�>���;�L�;���n�֔��?�k��÷�='V^�k�Gjn���v�K�7�ѦOV8�G};��Lqב� L���)��W޿xY�E�������n	�+�� ���%i���uw��Z�3;I:�͉���ƨ��������>�(�{uZSeP��lUlU+�ijd�����^�˧R�u���(�[�8A�_��'1B�x^��YY�FsFXG�%�a�Xo�a�2��ƅo�S����J.[��\�6������x rdZ?�h�Ћ	�I[����(Z�/jel���54<ov�_he�n�48�"�Y�U�.9��黦57��� �����f.]ѐ�]�n��'Jg���s��U�y=ۀ�\�۷a_~y��� ٪ �O���5?�I��H�vҋ_�cY�:�.��л�c�:���ù�c�nE��]��<�$S�T!��6�^Md�Pe�u_d���AL�����NS���8^��Kg�4����ox�Ah����"��[+U&� �%�����R�!�Ijֈ�ѫ���4�'�����u��$^�핿9\ъ���Fx"�US��+���"^�C�TIp:��1�ۑ/Y5**���02D���𾼹��,�DƟ�츱j����J�H���#V�gH��3Js��W8#V���_&������w*R$��]�M؅lA�Qm _��9d+�c��ʡ���P9	�F��*l����m�٩����ƶl'rc�9�H�~ڿ���m�����r���ƺa�����Gߞ���� X��I�-��� �eo�%$�.U�A-�.b2� ��E�
(�L��I,Wz��[X�v�|�w�j�/�s��`bǀ��H| z,L��ʌh��+�ҁ� U��V�����̱&GɭX��ܡ־Kb����R?vy��6f��E��.�>A�zq��4��<"Ks5�u�Ik�{�� |�H.�)����@�=�_��È��)Σ�{��� ?�a�z�X�:�U�fږ��/�@�N�T�F\[yo�<��ø�U�K�8&'�p&�Z�/b�ɰ����.�G9k�������|<p��]Z��/���4����
��z�	�\�wx<�����,����B��{����2�G	��pN|��T$ZV��\����g�q�{�Z���^ǭh��r���-��h�Ǟ5��=�"?q��Io�6�`�/�1������V�J�<�+�9���d��w��n�87��s�	G�JE����\��N�T���/����a���ɜ6��=b(a�q�,i2�!��1ӦIi�y6�r�9��EC_�Y�q@k�Qm�C�=��ΕKf�%L��t��^�pGW/�	�XkM�&+K��H��o|\{@�%"v^fI�5X��}}F��<�I�w��	B�ɠ�%1+꼰�����ڙ��t���*� ��ĸ��c7Ϻ_��-#�N���R�Q�Q�W�q%�������I]�mc���Z}ٻ/fD]�ǳb��E0	�'��|�*��e�������;f��K�lJx]2^�rR�� Ǻa�����8���=�z�C�H���6��g�^�H�9A\RҎ���=r��y���$R'q�_m��^�g���U?,HK���,^'ˉ�t�����;~g�(ql+����h(��[�Al ��j�t�<n�3.�ֺ�{��?�/��A�Z�&��S�����ɩ��?��˰h�H'w�6"�|��(XX��?��R?�����m�_,|U��<+F6��(�^�Mf�a���Yi����Rc�Ѻ��{@�YHǔ�Ɠf��G_P$�ڂ��Z�6��s4�3L�T������z�D��]!x��`����i�j�JF��;�Ƨ�n��M�y�6��d�����,��{2�o��%�"	�U��6L	-�H��g�YƐ�g1��g��u����CL�$��]�� �"�M*��ѥ"�&���^��`�*�E]��,"L�/,8.�7Y{��bC���&O3^���Js�~~RD�txec�7>=�<B��k�5�B�`�9Lқ��D/|��_���h���W~��t�<b� V����Z�b$���k�K$��$��9R��\��XS�V���c0�D=hp�Bh=��6�<X������l����N�.�,vR~�3+�VŪ,X�V�3&���Z��� ��RN.���d�
�!=_�|��SƟ�I����=��u�0$y��z:&�جQ��>%\Y3��ҁ'g� y��N�-�KAo��+�S%�T�� �A�ٚus�7<H`��.��Sf6E�3`�
�6d�~-��n5�`�{�����W�QQ�E���#[����-({��0=��	�p^̧��/�Ӻ9;t�^�Sk3s���5AX���`�$tY�߾�S����� VN���@��@	�!2�n��c�����e�&���p�w2����o����ln�1S�BK���y�m(�4i���� )@�|A�A7̽H�����繭��m��w��Z��-�b�c"���|<4�C�Z��g���fE��o-�?�ZG"�)^�<�4)Yӵ��|������oʆst����: 8I�^�
���||P!�YX�)�n�ָdz7�X�I���b�	Ěy��#��$���_ɻj����jA�50�0��%�R#�<Ҩ 9u��4&ʅ�'5>
7�0k�vU��@º:"!yfߊ�[�k�3��r$������0MΉ"i���cX�6ߊ`���t��n�2;������*�׃���E�)��h$S����pre���,|_��^Gv�^�UN
�>Tzҟ�!*��Й�$C̃�vf�q[��&�>Pn#[�7Pg�o�s��"�9
�Y�j���4�����&�e-妜+��J$��<�*�L���a�+�mӌv(e@�b*P�7���6>�?@- �*2.��W$)��
"L��Um�?��DX\ϑ��д���گ$IL�1��PǷ���v���Ǧ_}�7��1�f^W�7랸�j⠿�j����ΦC�ϋ�ø����#� ��ݡ^F��K�/x�E�/G���b�7} ��O%�R<��Ԍ��D�Z�	;����}���:�4�譊�b?V��Q�(	�ZG��5�lI�p�u���W��ҫѧF�2��~�O-8�����H Bj�1��<�YE3FL�`%;����o&ˁ&a[���S�h�ҾNE[�L�\BDw�C��� f�4?�nHh�f,	#��[�� �Kj4�#ڇl���5(y�v��hY�o���b�t�Y\��"]t�]^5+�?��#,��v�"���W��bi�'����p2sa�I��=Oq�P�U��aS
Ƞ%)?�t���SQC=���B��=�5�YZcv�ˤ�w�F�GF.���}�:Fí7��H��vzJ�[��ˈ��������/qWy7�^RH:�ߑ�'���]����ЈK���b�t��2��*�-�nC��H(?b_�o��tn�izw�ϝ�!`*��u<�R4�у4�H$��;
w��4|�>���DT�RQ/�j�*��)~���k4��7�!W?@��Qa���`q#��c�ǄL+�C�,�$޽���|�=�pY��[�8� ?��w'+��A��x}
�A<���k�FF(�8(�(]2
6��v�)y&���s�����ʙ`H�.��o��ߥh0`D�E��,�4��YބC�}��b<��߲`��1�|DpV�I�_�\z9  쁞/���~pj[]�>F�O�x����p������X�
�L���㔥�MFq�-/�*Ƭ���m���ƕ��g7}�l'��p�5��.eA�2���tL�8�$Q��;��.λ!�/��A7�"T}����#Evo˛f�G�e�Dr�6���xܵ(ԑG�;)B�ǲ��m�N,x܆���86�%S(T�Mb4F���e���CO/c��!�{����k�Q�ƏG���_�P ��C� �53��`3HE�܉����������!���`�8ѩ�z�j}4��C;��� �nn?^M��6'\��=F�s9�3`{��,��<��=��QN�6��o�YH\g�R��`�1�Д�fZ��տKV� ��]n��m��ɇ���!"1�#���f,�&�]B�"H�d/�Q�.['7���^��N��O/���t�[�z�CD	J�e�7�a<�ʉ����>NaS<aҗ#�D��� ��OI%��GD�d��8Ar�KV�*�����b |v�g&�GP��^���59ѰA����"�Ҥ��|���;p᪦=k-B�8��œ������*w�ʢ �ЪR��3'CD�&��a����F�r��Vٕ aYR������dj���-��D���@,�#�ߤ����J�0py0H:"ZS���Q�"%>���/�N�g�_Uy7�,�)ٿK�$��̐S��cT�A���������78��`z�[�*�S����/0,��\xd���-) n1�`x?Ѕ�����"�Q�Q"���B���-����,��&��l,�H�O�+FT���p6��*�k/Y9X�:5=���˸���Y��O�}��x/��I����b�[��On	\$�:��l��&�A���C2�6�J�߼���n5��S�-q�]�uȑ�i�v�s)e@�y̹o��.�����w��s�xZM�X�^B�"q�)x�h���Z��gԉfA*:o��U�
"�]�8X4��ӱ�|'�����oF�ot�d�a�  4I;��
�(|�EW!�R8���{���4��7�o�I�T�^����ʚu4�#d�$�r��HCN�f	�\�=��0r��!�#u�j�ټu#4"YX���9>uv0�p�gֶ���A�'U|O�#���eN�D��������E�pFW��-����\��\�S~̓�����pP����#��A�d�,�j��$��� )�]�x� [����8ml�VQ�^���N�`+�l��O�b!'��s��LV�^M;���hV�ꇉк���Q�cT�qL(�7��)S�Ό�}�LC��E��Cw�ռ��B�z�����
�{��V�}���B�zOB��N�Ww�j�D6�
�uvo�='���pU�d�),���W|\
����L��L��1%Ǜ�d���	5��10o��
˾�gf\1d�v�S����D�"���;L�U��-��1��Q�C��0K��LB������G����/�XIZ�V�KO�/�;�%���\��t%R��fy�(X��o}�V`�R1I<~Ѳ lד�H�%Eߡ��$����`�
����AE�'���0��J�I��aNcgs��u-S5��V�QwK��-0���f�y�m������}	(mftO�����uny4���Y*������@zf��K(ՠx������+�0�ra+˳� W8�s/m��sU܍'*=�������o�iq`R�4��9CD��������>RW_��R^�~#g�zi�2�\���J,�%e˹�t.IK��˼g뾁l[���$K��!�A�.�_kt ��Q��V�7��ow/L�aA�_͆V�q�+o�Kp����������U�x����h��6�(�2��o�B�eʠ�rm8��,���l�6�s�(�hoM��T���������^cʹ:�/j��1c��ي���[�w�PT���=��N蔣R�3|{8�=�ە��t�&�4�!���`F֩�.uj�^#�������n"��M�%K6���$?O�Кb��Q�{b�>�6��RȄ�f�6O��9�H��;g'�%�O��1$@u�ûH7�X�s�0�T��]"��Ps�}T��2AH"���^�#��Z�]���"|�]/\��.H�G7�!������Oc��(������D��ceH3�7n�<8�X���:�r
�"���D_6��J_+�o]��#����{�l��&��V� ��D~bT����(�{ I����i楰��(�����͙HÌ�t�Ppo]=x��lPv�G�#j���%?6�~$r鵈,R�œ3[���Zۊ6?�c��<�Q�
�W AZR~,ǷK�diQaQ���S�$Dҟ�?F�Η����0C�y�:t:V��6��Qe>U��c��~g%�ey�lK�]g�Kqy�� |�SU"�T�ɛF}@�	�H�
7l3v`.��	tS�� �c�0�:_d�-ݟ�ne��`,|N��^�\�Q��)��%8��8E-X��`Q	�ڣ��������_��im��w�̃��kc�6��5qhe��=� �Y�A:��P��1�آP��~�V�CX ���Q>�n�.v�McD� D�&@%}����2<\��幼��n��
SK]���̟6A��E�[i�ջ'��@"��3�퀄������K�+���Z�Z�W��j�"%���0�E�pZ�6g�<,fu�)o]�4��&�"�{��lQU4Y����$�|��ʝ-@0o��ctK���	 4 �I�,~
�'L|5��!蹇HE�^��7�PI�䨎�ڽ@S?����#�g$�je��A>�����Mؠq�10ͪ>�Ua#)ԨP�Lu���4V"��W��>:[�0�9 U���0�!�";��uk��1�����d#�VιB��.�X�"����;�F���A�;�I���Zk}׳MV�1a)ɭ�hT;���Sr����\����ޅv��U~Vz>�L���9�����T'փO8a���������>�p�#��PK��o3v�ļ9:�r��p���z�,%��.��e=����o��z�ؽ�L�*D]�/�t�[��Ӽcepm�*�x87�6n_9?ps;�Z>��ˀ%WM��TS�:�)Lʳ8m��W?�?tD������M��}����L�[�g���}8�����oVg�,a�^�����B�jq�����IƦs�������6�5Wm ,dF��{�Wx��AE�Cw�)͒�2ϛ� ʌ�%�����%A'Z��;�l�ͭ���j��ȩ���X�!�B(9�Zw��e ly��:/����<��v3ܬN�Z��8����v	B��@����Yu�F|��%kl�  oO~,�V���)�S����>�[C�\r fׅQ�z �{�?�hA�	S��[����{Vt�SL�l/��5X7PvA_h��z����F�vY����R�X��F�5[�������@'��C.`��Sn;d'�
���+sOEyR=!���l�5�a���Uqb�D��ggs���"s�m�����v���ק��ŕ.<�F�H�:; g��M!�xfSv���[��Y��S��>�J��q���Îa�Hj�$	�Wz������#�иu�Չ8b���b�*���Kc�x6�b�b�o�کn+
[w�u��E��*�F��<�p����x�ߥk��w���|+�P��f26�Q2�n_�G�Z�l)����q�����Q�9?p0wQ�����ė#�V����+'z	,�A���ì���'�%�\8��+��+�Tð�I&}:��<��3i�Fv�@8X�]b���	�)��Q�	�Ws`���Tj�^{֟tS��.�`tf�����N�l��<�C$������V��VB�A��1ھ�p�n+��eozitd�x����~��i]yF���b���.��f�,c`
$���g����F�R+��XΣnw��)X�A@�`�ay����{1����mHP��8�X�g���^��2���_�����0�XRm��2tN�?VC>���GG�������_'Ffo1���3T��u�F�G<�L��-�3�F !]���� Ty9,��ū���ń���X�QP�!��7f`*�ۈ<r�xC�	���+����ғ]��k�g�I���JB�����ro?�պ%M�;�q����@hk�x��-����ջ��[�b��Co���p������q����(u�0!w�b`�	�o{<t����I��[��9ׯ�鴾����@w�����6J���o�a��rN�B�-ci/��wi�R��=���P�[������c��d�XFX�<�]�(y�G��pȒ&�Hc��U�	�\��tY��=��~��p�!���:��Pa���v�?�A=NQ�G�ut|1���*�l����3��'1�/�N�~0�(�qB��2s�<���IJ9W6�<{��Q_�zq�������C���³�TKg?�L3�3��&��xZ���>/y��X�9�pdK ��,Iӝ"�\��%��f�@iXPռ}^�OꉎI-4��൓*?z%����]k��v�������u�Ȁ��A�1{�^�9��cؚ' �-�����Q"�	��e��_F@�=oQ
Ϊ�N�����`}� �f�F �t��mk��ѫ��*��A���P��zuf)MPKYORx�`b�Q$����a�. ���Q8�z~�Ĥp9�x�=�lw��ܕ��IRӆG��5�UK��w��S�Rȑ�_.��^`�1g�}E�v��m�� 2,�(8�*�t�d앐Y�g��lL�й5ǭ�R��A��Bx��t��
â]�!��(&R΀m/}�A<�6���IO��?��eL�{��q<�����;��G>(Q�� яSl���S[mI�,�����S6_e�(_�RMG񛺌@��&^��c�;%��2������U���t.�Hn�PE������r��ۚ3�.l��2������E���8�!�^�`C
9��x0j"�G܈�q����n��MǊ�6�	>�U��!�'�Y�{��s���d�#kԄv,j6`2�j�9H	o;g�$����1����H(�	Մ���(Y]s_T����z)��Q"�[:����+�Fˋ+$]�"��o/�4.��A7Z0M����� �O���y�l�|uDN&�e�Lh7?c�<)(B��SMȣ�mXx��<��D�^��������ӵ��ɞ�����%wP�V\�N�Bn�b�����l,#13�����F,�ς����Й�?��E��p��=0�����?Ř�����-Q��3�Oxt�VyR�Qz3����+/���q3���g��?ן�c� 2<JR�9��|�\do�� ��=߻��#@��p��'k�F�0t��y5�F:�!��$oQ�L>&��T��ggV�Oy<�s��h�K�/ʱ��S&z�T�\W�:e���7� `����L SgU5�T_إKp�d&Nn-.9nֻ�`����l���X6mQ�Չ�·����-�#g���C�kֈ�Qxͨ�P��z�����ԭWk�<��� 5")�Iv��7Y�����f��c���0!�r��æ�#�Bun�C��~]�q�+&�l��1)t2�#o���)���jn�f�SK��3���iE����i�����L@���J`�zߕ3�ֈ�Iȼ/��X�lZ�5ù�ğ"6{n�>F���9Zl!dgSu�f&��o.�'���#"֔ˇ��64�F��V�|l!��ޫ�o˞�t<�Z�&�{ e�eI@��
,��|��W!�FJ@Y����1�7ξIĎh=ю��Z=8#�$�H�������螼��$�0^�6�0#��ͨA{uҲ�4��M��8�>���0,wU��»�!���<|k-����v�ϪI��jS���X�#���D��G���hn;I[����ׄ�W�"�F)�M�h���m�vr�U���4��1�v��Uo�>�my�}��,�������y�W���r�g���o>��#��P��o��ƘU�y9�Fk�6�e�=H�_$4e�֎�=r�$޽��*y�� pf�l�
��Dfe�YZ*��7r�!66�?A s�K���ܥ�W~�h��F���L[��m��t?�-0Dy@.��u��
�s��P1�L����1���ˬ)��զ��N��)�1�^��L�_��jê��k)��̳����-��ڸ	��צQ� ����?���L@�xE�!�����]?@w3 [��%������f�m�Z06 ;Y/���E������]�C<u����(*�XZ�☿���l��%~�T�z��ճ���G�6�?����G8��k+B+����Y&�*FM=K%\�(Mo�M聧tƚf�SO`ҟ>y[�8w\c�f�3h��g ��?1ch���	��[�6{�lgڭd{�l`�5�n@v��Vh.V�jN�BdY}Yb�c�����5��l�5��QGw���l�x&£l�'^��_H�s�(Y
gT=0��Q�Iviza�����e��<��5,�*���ǜ�>���z��v1w�خe�G.�����:���îɱ�i\�v�`�[-�Έ4�o�+����G�q8�T�_H[G� Y_ԈQ��ި�ޔ!��I˭���_b���SՊ*����8�ɴ|b �oh1Gn�2�w����6��*/�ޏǳ<e���r�	�$�w�|U�Ug�nQ�������^)_ 4�2z�[6�b��?���Q�v��/��#~ܜ��@�+�{L,�W���ʚ�݇���C��.8�u��܄s+������}K�<!BP��.F�8�M�]h-�ڐ�)��(��sOZ�W��:���pc�PcGߦ�	`e�P�*��k*��>C�t�xj�yb߳\��2P�1�|$p��)���=z���Bק���~q��]��F._�كG�'vc�!�ʋ���
��ѓ����B�F�`+��ZX�ywp%����A�,�2B���,�漏�).�m�y������Ue�r2d�ܑP�������?\�mT[�2�"X?�">57�GDj�$���K_X��|J�'�TX4�uERG�L��ܙ>xB�wT!�	��T��T
�0�W�<�m��u�]�i-��7a!ݞ�f���l��rq�t������}���`��/t��G�ߺ?R���u8��C�����M����������x��-|O;�]ek�v�Mb���C�i ��9��	T�Np���N��E?0b0bqhǠ�ct�*�����݁�2����������@�����J?���A�Oa|CNd�y-T";w�F���X�Vc[����}�`ct�Od�fKi����dS(��Gu��pY��jGocū��t��m��t�xX=�=~~�pgv��X���Ѫa�z��欫p"R=����8�&p�NI�K�����ʼ�/Y�[��Ρ{�~Q$gxWE.�N�V�"i5�D�H�S�񙲙��$�+������4~0.��"QK���6������B�-!�}���~lZ�c�ӐG�������B�y���˶��P�^iYW[��<�y�搥@��΀���j�����g2Ȱ.�&��s�j�N�wmE�v���� �E2x1���ID�I�~|���2b�J������V��ZvY��Y��~d�f� 3l1���`h�B@G�PY�Q��K��+R���i 3���4��e��WJ�߰��4�	:.�@�Z��3[��!s����D�0�OlcNS�@�,/ea���v1��ƚ�l{a�Y������$���&i)�=�,hݘ˚�+j������mK�q��5� �u#�ҧ��2�j9��x�](�C?
���Z�֙�ݠ���e�,ON��
���o�`�n�Z���xC	��g���WN�R{30�`�4eD���*�I�����\=  W��aҬ�e�u�H�����/+͍��:����ph
��-け�u�8G:ɰ&GL��F;ΖO߻FЫ�&?�$g"&�������\E��}�<1O\N�T�v�oz��ɜ�)A\j�HA�\�nn��bz�-�<�"��\�")���n ��i�xz�:��]h���ț���_/z��5�ʱ�%+PĈ��FU�*��V��IN_htQ�x�5*����5��ej���K8 �t�2�=���o���ŷ�N8�)jJ�Ϛ�_|Pd#����A��?�$�U6�^J	cF\H*�Z���Rc�T���i�B�Vk�45<�B�Pq�ͣ�M�H��`c��6�KR�klS_���9!9j0��wO���xgm��"k�Ԣ�l���f�u|���Eoj�:(�x����6�s
f�i����u~��jE�c�
�0P�p�b r���*g���w7��n�Ea�h^�,�Q6M���P$�Tiq�Z������#��P�,���ц����q���}4�I[��\!����>u���x8)J���<�_ԹE`�t�k�R�J�K��;�Ջ�T����X�G%�e��,�r�V��|sy�3Z���6ro������:y�������r�+�b�!~�чc;��2:�����XL��7�zq���Ƶh���JԌ��Uٙv�;�a��"���؋9�5�&~��W��sO�0�aH�m�W3�����;�!�<���_�їL h��Ι�H����X��;�!�y�;�zL%�2
�bV/��H33�m������K9j�?��U�cpe��>ڒ��IǕ�����H+pE����_�X���!S�����A�%ی��S�"��A���J@ɖ��R�!��?��_�-��F�m��V08Y�����u�����G�F�)����1��`jV���;R�h�����TsTQ�:룐~(��7�V����}���QPf���[��b�B��`����
��D��}JwB��QO��NN1�W����C�y
�V�o܎gƐ��}�d"bM�QW��m\	�"���C�-1Ċ��,@d��	t� �P�������J�&�1�yvl��W���v��"��{�G�!�B$Z���d�uL�빱�p��F3H]t�f�"�d�U&�!���=��w�+b:	|�r##bSt��궪���h���4ؿ���@�O\r�ׄ�A�{s?#R����������s��_I���wP����a��ZwIX�{�q�;#^b�P=��&�J��Ǚ���ޞ�$k�u��	�s��t��C&;g����8`F�W��E����!�s����Tk�O�2��ZM����
-�����.���q�o��p����MU-���i�
r�'��2��g�ھЎ?�Ea�P�$��4��U�͇'^�,&�EyG�ɸ��voo�1�4�w������㈾��y�R؊�?�~��FA��Ţ�R�ϝ���-�I��͵ss�g�=�)�W�� �ʎ>�4�;`�"�-��z�f�D�~��X��萍��;z.Yu�cS�B�6#E�F�z\cɇG����r������:B�1§%� T65��f�\���Ƚv��g6ϔ\`��J�@ ��i�״*\2X���AQ��.�A��P��=�W�W~i��t�S�;%5��2��CŚ�DPP��q��۳\���'RtP�/�����C��X���l�VX�T�7��O�^;��P��bu�����A:�̪��;�U�� 
7�&��^6�����;��x�U�e����;T>[�~��*%cf��੆�CTI�ɢ���q�ٹ���Q��X�%aQ�6�Cuo/^�濧�Ѹ��+n����"�?��d���B�^�PCd�JpH�i�������Y��B�'n�0 �����'�m�Z��ƍ��_[��Y$GJ���h�ў���Ձ���JaZ�W���V>�_='���k�a\�w�Ej$�y�;�l�9���t_��1d5j���v�=��97�7� �6l9P9j�[�h��m=�dY'���9�m"~Ȋh4
@�%���q�$��h1諄���uR���u� �N�����/��ej$0��o��.P� o�JEVe��z6�7��zTG�[ƎL��	�>��Xƾ�HǮ��Hj��z�e��^|i��._+�պ�ε����j�#��̟����X���jBb{�� n�y�JfIbEܒ.�C�����-��*A�s㌦���{�ڃ|�.��%��@��_��?�H�)<��{��5 -{��(|���rU������Ȉ�>��y�tؤy]���GMC�&S�U/�&o�'Ez�&P�/��+�x���<�G�.S��)��;�<��]ȼ�/�̞4��p���O�.��	Bx��e�<8P�B�H��S����K�J��˫	ٶPN��_��#Z�i�����6}��O{�8� �Ǜ��OCߑ0
��[��h��5�1��:R��o�$mn�݈g�Q��[7��J�P�+�������f����>������J���_�!\��'�BY��ݧ��t r�&�ݜ������!(�_�q��2��K�ߩ�I�B@6�	]�f��_)��qn�Զ?4bC��n�@	�K�W�L ���"�k���6./��jX�ݜ���@KM݊���ޝ���\�(%P�f7z/X=8J}뜉�`�I�Ke�~��7~�%C�&ꪡ��c���H~&��m̀�~b���������\gc%����-�7��Ϡ
�WQ�8 ��}�!���������cܞ�/}Ǐ�f��!���s�t�����*-|2�(X���ef��AKf�tx��ʗ`{���eai ���8����$ı`0�%�ι�n��m��#R �g�p;���k��$� 9�R��_�^�V�g�ZE�C���F j,���w:t�����g�Dl�Թ��1�_��A�����t~��P����>������'�/���A�J?�!���bw��9�u}�y�W���D��͜�j_�(sɭ0������ʆm�A&,�Ld�j�6�zN(LGIMԍj��n�WF�u��cW��-�/����BV���b�uy�P��u��(J�����3:>�ܻ+1� _�rzj��%�!&�`P�ө��jo���ud��4Pln }�M���6Y�֗b����9��b{���U\Z�P|�C6��w�nH�_g�*Ԑͭ/1b�-����C���l���~] �3�������p#h"�2�������˘��]˾�":��/���.��L7�i��P���XO��$�&���lymD;��e��T7ly<�b��hȰ���=҉�Dݢh�[u��浢';�4Bv���F$OV��)�/O&b�	f�b��9������/ΰ�JZ��}�^��{�rc�p�.s=�/������E0��:�l�}L�|��s&�R,h3��s����_t��Ɩz��ˁ ���R�`��|\d4��n�*4�b��Y�����|I�0�M�y�#�:���QMJM>S��!���#�gc�Gy�sq�N�K�7h�>
�SSx\T����J��G ��/c7*�>`�#���S�0��!�)���#d3�-��Gn#�L`�v���r��Q����//ʛ	r-V*R�ҏ�X<P�ޛ��=W�ZG��^�́k!�� �5�n���S���YP����E��/$�.�_���^�s��� n;�ϋ�v��x&�?��f2[������vL�ngR�SX�U���۟�9��Þ�i� �%�f@�9DS!�+������Ք	ȩ�g���TZ���Pp�"����0�C�]Z��g@��f��yo[b��
�"C�a���4W��ӣ�O|Y��kz�o�>�t	{��0 r)�I�}A
y�y|��!&R�F�$�m:2�f�O7$�MI�S4�P)��yb��'#i�$����zwl�����Ke2/��0Kogѓ�]#'�?�!4u?i~4�e��U>�>�eT0�UB|���*n!g\����k:]��{���Ltϗ���R��,��X�:����E˜�(�;���I-���ױ����V�)G[h�����irSQ����a�:��v�8tU<*q>�l�,���2��l����@@����sT�>�Y#���PI��oٓʘB5�9x:b�� ��pmݪ��l�e;
���Ϙ���3*B�ԉ����������en�l*>�7_c6���?n?�����ID�W�*vR�����LH�m4,C?�)�DF�Q�j1P�"3���(ڝ�HLr|��gV����z��oi���_��^Eb��L�&jP�v��&��/�񙜋)5(�� ����
 ��>���y�dx���E����B_͐��� HW�%K�.�m����KZ�e�@7EӔ2����L,R� k�E�'�5�I<���:Y�R�.�<�0��USI��nj���%�<�Wn������+iW&��<�k��2HI'���漣�n4R.S������՟�B���i�D���@��Б̘�A��Lւ�����3��]�Z�>��}�3"p��WEb�Pg�Zf��g���f��Ao��L��[�"NćmF4d6��Pז|��G�X9Mo��t6��`�N ߖ�I���
&�| 1�!�tӖИ���H�
>�Z����~��wG�à�8�Hg >�5J��f��\�_��	'Ƥ�.a��[���R��Ci�PO(�&�q�'j2������I^5(6��P���|[_0k�qUHl���C9�i�ǒK�CLG���I��e���/�1�Xn�y��K�A�@B[����\�5%7@�f���X��}rT��	�IA㲥O�>�K%*@��q�K�
���̾�	�n�,�H��g���*���Hc�����-~�67m{Q�b��o����QN�����b�6��}Jqf�p�(R��Z��6?�84�*���t�д��f��Km�xrU-�'�M�U�a��ǳ��8��x _ĸ�����΀�t���:�.-�Rg������w|����熹R���_�^t/�g;DS�(��t'.,s/�>�tS�a��q�gP=l`$ٹ����f��A�7���t%�׎����<g0�u/�t�A�}�۔��V� ^(��)Π(����d�����1��(��!�4e`炘��<�m���,�l��Q1H6s�V(�=YM[Yy� �j��5��}�c���������vƈU���,PY%���GK�/�����3*4�b�������٤����!Mf{`W^�~��j6��7���n��M�Û6�e�ir?��6Y�mjx{��K�܃=��%Ą�9Q6��~}H�S�g��.�t7�1��(W<�f������r]�����7��'b��x�"J�T��[b� �˟u]���"�/���.ߨ7�暸�! ��/O��!�y�3o D�{�eU|7�m2<=�x�@SOȷ���w�P�uD�V�v�h^ĵ��Ş[#\�����1VpWe��k�b��D'�1���I��L}���ϖ���1Y�ć�ټ�p�=�~X��+��,�y�*����K,Ê����?RS��3�(�ſ�"���q���h�l��o� F�%R#����d�~֋Ϭ�,���#��<U��|��=�0��yɽR:�Ӳ�[�8Q��I>��Mh���N�gj��y�ݾ��uK�����E�S�$dT���?�N�-���7�|5`SA���+S�S��h0ӥ�c�d:�a-�ann��B`QKͅ�o��Q�z~�V�#�G�-=�`��m�����e��aO�d�~�}���h~�k�D1C�56oD{�#�Yw�&��Hu�������Yv��9�{r=�V�anb�jϒ���Zi&������2�ê�cfټ��n��S_-����ϟ��E�j�i�0~���o@'�_k6�2�����֜���P�\�l��Zf�m��a�"ʺ��p��*oZ�(Hg�^f:�o�=m��R"j(󇱒P4>)�j��| _����o_��tP����w y��Iԫ�
@�	|Zbe!�

���0�֍m�7+|*I�x���Let��n�4#}��$6c֡m���~��2���{w0� =���#��H�U�Suf��4�7[�<Q�>�ժ0�1U��I�OYO!�W���s�kAF��������>+��~g9ד}<X�Ԋ5����E���)M;].h�? D�����6 �)n-h��ڱ�rF�䁀���vN�U�*�>)�s�3#��  ��u�tW�k�������>%�#�;NP0��o�6͘�0J9����������#�sre"窦Q(���@��:N*��ۉ4��� ʝ�g_eU�w*�g7�*63B�?ծ�_�6�p)?W��9my���L�&�m�a�?BuD�u��M��)����dЬLTr�E4��_�!��#Ԧ4�.�eF�'^8��_j�2����}���<�$��07����׺�	 Q��S�u��axX}E�~��(4�wf�T�� �SB%�.��r/��*�Z�];2s5͒P���=��W@b��q�(>��Z^���~�l^z|����������ہ۬SD�$��8*Ĵ��o#B� }�Y:~�F�k%p���p�o��B�;��Ʈ�S�-}ҳ��[i��\w�f|�b� x� {��?EB�h(�m	3,[2������F`lt��5=o�vƳ*h����~v9��l.Y��q��΂��
�5@ܱ�I���d�\�e���w�7�!'3DV����s������=Dud����a(�᠚��)9b�I������k���t���jv�L���<�Q�.��ڻBa�: ^�BD��})vOЂ[A7Ո�EB�?� �oa�qL�%���Ho���HԜ���r��ި,���8����ubU��gJ�*�����ȝ]b��o��]n�&�w9+��J�Z*�O�+�f<�pۆd���(�0�3w^��|0rrɛކ{��Q|��[��O�)s��4Qj�L*���I?��Qv�ޖC�#�V����+��k,��ޒ2a�����FB�� 8'����ȍ+%^r���}ߟL<5pV��F��V8}�U]'��n�Z)��%��ɹsc\��_��N��׃*t�dOo�:b/`y$��L���AҤn��C��i�xw��n�Gu�Fe14p˘ �t��z�C-��8��� ~��]�F����ṻ�,�5뻋Qx�
�Vd�EZŔ��xFFr�+KX�@tw�+r�NAiN�� G�v�zpԤ=T�m-����᠌�A�#�p2��F�d`��1���SVWm�m2��?{W�>IG����]��)w�_l�TQ�;��T�9�uY��G��L����'�؋�!B�O�hVT��C�kH��F|�ŉٯ��0����!q��f�"�� �.r��w�n'L�0rٮi/3��y��PԆ��2�沓��l��t���l�M�.��AղpR����-�W��oU��Byb%�wC�[w�UI���O����*�����0&�!boǴ�et�i�>s��;�ݕ��j�m����Xa@�?�] JSj4��+�a��N���-h�Z��w��w�����jQ�[ ��ڑ�c�d��	����m(^��G��rp���~sDcYZ��µz�t��M=���~���p�Ù�l��[��a!4�ʈ�q���=3������b[��H;�P��/m���nO�{�`$�m8EB�N�IK*۬i�f�\Q�,�I���$}u�$�z�퐕�d$~�!��6�s�+6��ï3�B~v�f�-��~ �c?���Gȯ�G�d4 y��JQP��������$v��椈6�Z3����j4��'� 2\���.���j�fw��v����,� ��2Gd����D�^\�^�* ��^��ME�� L��l�-mbYJ�zx.܌�t�1)d4���t���O.�G/U�Y1r��_+��C���63��4�eN�s�F�����gN5@L��]3��)�5�a�H9YD�6��4�N'.@*jseu��}��1��N����{u�>v#���߸!��:-����9h񱁚7g��-�H�I7$K�� �ɷ���fB��F��9��x��O��"���j���I#���Re��NKȐ��.���x#�ꊓa�WY�t�ќ�UNW�%3D2�`&�{X�e���I��؛}� 4����c�u(	����ie�͡o�:7�����QS|\�c�ukM�:�W.G�y�FO�$Os��п��Գg6�&_yƳ�y\��P}��sO��T�[-�����)�n�\�9\���q�Ir�AA1���/p�))�ȑn7���?�z#nξq�涪����l���tk�籯1��޾���UO���L���g|?P��5>��`���<jv֔K&8��c�'�ӯw���J<��˛8��j�/�Ϯ�z|�đ�5@�X�S_ȷ����#;�	�ŽH>Y�B�MRw�
�z�i֞
V��$5Pt.�$��@��n��&cM$��_�:k��`lg�n�5S�01�c�6��T��0͒��Ga̵N_u5-��Y��nw�hQ�}���1#�[ǯ��}�coF}d>q.$(��q"(E�6GPJ�p��%j�c�!��϶z�(��t�p=��h~Yz�p�<���-���ah?�ʯR#���=.�eN�aA��AF����I�w�/t���U`{w?�$�T2E�E�vYq��i�HY�c;���ղt�$$�ɫ�۶����t$~�:��=���6t�]�V��B�g��x���t�D~'�c�Đ�=�z�:�@jyi��˱�9P�nz���l�����kx�ץ�?Yj��A�n��2�^�̋7�g|Tj_f�w�X/vB��n ډL23<	��)D�9�Y?���Pέ�Ǡ�;�G�ѓ�t�Y1��?=q�;\�1�@H}���[�v��G6�Y;Z�&��+V����%3���4���1������'l�f@�Z�=�3U��|T@�o
D�,���N��	@�vme����p1����Ƨ�{|�h%$���1�_���e��8D�h8(^�^�N�4��0�[K�6M�p2�r���`썹X9�6x�n����y������$�e���e��Nru˯��B���I�w��I9�V؛�X��1��N~n�3K��`+�a��J�I�q��� {���:۬��u�Ķ�(^��N�(�:�&����2z�b���uRŏ:�̀G��`F�L�O���&��]�g=zF�z�n�M\���}n&xOWk�TD3��*�:���)�~��#�R\���	�^�J�͈o�݆�w��)s%�n�0���r�z���57�z���H>������癷��ݱ6P�&�Ո��UvL�VD��Q�C�W�F�5�{���w"H�j�r�K-#�������ZN��߮Z�Q��Z8E#�j�ϵ��|�������%|��B	�P]�j�	��HE�q�)�|R> �!�Ni]Vfk�5��
�e6�y��(��ݞcc������k�6�l�s��`�<��0�]O���xIl�[Rrk�����!�
|�$�E�����x߶����
a�i����04�-'E�s5
�P�&�,O�3m����eҀ5I7�Bh���6�C)�,�w�M������$iq��Q� �I=����,���!SN���ޝi0���wO����>P��˳t�J�߹�7���\S��U�k�k-����ޚ8��"��n���\X��%=�}�G�A�W��n�nN�<rj���i�:4���v"�z��r�M-�.�~�ָ�^ө��:l�����L&Ű�U>?�N/��v����E����T�1V��aTt�"�[�@KX9VZ&yAbE ��O���a�k0�2A63�Ĳ��;�&<����k�W��2I �5�gbH����@>;��1��e����L@S����V
o?Hn�Xm:j��r9�P8����~�2h���m��fH��￢p�W_���u�x&����S�j���   �   ލp�F˸�$�R=�1�#l����O�ToڬrN�'|W�DC�O���]�e�����:Vؽ�Da�w5,Qlڿ�M�F�ilZ���T/f�l����!��TI\&�L	���I!����һi7&�����o�x��f��T8���,O���bM�HR��V��x�Il���>yUJ^2_�Y�C�b|ެTf!m�04Jܴ�M���F}�*�K�	_�ts�\`�D97K�p��T��B�	5?��0�)Ҿ����6`�C�I�m�̵9��]�c�B�L���C䉹|�z���#CR����_8D��C����$h��ѻZ�\�)�Y E�C�I0<ĆDY�*]0�|9�)ˀm�2B�	�V� 4C�l��,ŌD3��!��B�IY �z�ꊘT�\h!���1ݰB�ɯ>�h$3�Ꚋ7��H��ZLB�I���I(�JX�t����`���C�ɖI��D`�YU��=��@ax���>	$EJ�AF�s��ʻN���QD����O4��V�d�27M>}b�ǚ�ug�O�� �J�-D�.ez�,/2�\�@��d��O��L�\�4ᐛ,5�șv薹���AC�>Q�1�S�#<Q4��-}���"��990m�g�<QP�I 2  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   5    މ04�̐��%�R(O5f��p��'l����I�l���   ��@ӌC�A+,ɘ�I'\	~�`%Ϲ>   �   ލp�F˸�$�B��>�1�#l����
�޴Y�:��O��d�����	�����"fŰu�pph��^�wS,�ش>G�6$}�8����
x��ј�R&?&����[���x`&�j�"<�C~�����Y,~(��v��e��W���%���36ڱ�-)?aQ�E��7Xp}BJ�8���D�5{>���N�!��X�Ӻi]�V�Ϟ������ē��.�-!�ph���Ȯ.��x�ȓ�V@".V�>��`���G@�ȓ]d|z�	�i.j�i$e��N9�ȓQ��
��p�GCO�kk�����ZG�<��"��(VX��N½,�V=�eH�<! ��/q��̂0�� n��iI@�<�P��i��`���?��%b���P�<��*�=E�2�:C�"�D@�0b�M�<���c�P�Cc٧o58L�1%Np�<I�"ϧ3��m��->n�a!��o�<���f���'$«h#�+WfD��h�'��Ň �¸��O�=y\������I"Qf�n�󦹤O��7����rX$��N�1^n��6bD�_��➀��I0��B �3b�F�d���
q�9�'t�Ex�}�'�R�j���2������6�|���'�L�k@ ��<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&�   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ����Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�   �  �  �    B$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�U曞@�VM�P������@��P_`���'4r�'d�|J?��f�s^hy�&A�x������ b�8�`XTv�|2���,�
�*��ڹz7"a��iRȖ:[�Fi��	�[ڀ3�F�\l����S�
��0ɂ��O��d�O:�d�<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&��|�����$��::�i�V�%C���e�Ԋ!�lK��O4�$�O��d9��~r"&F�L����� �45`� ��A%h�d��o�&=���1���Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�Y�P�{ � T�>�@� D�(1! " ��Eɵk��<�s�j �M{��$�~��A�(���4 ��7�*��2��y>���=���O>˓ I��"��ߣo��u�)9?Ԡ��F��r����y � ыU6��ȓ~�p�k%��^��1� �
$F��ȓN�� ��啦 jN=H�Aއl�І������(����� #zy�q��K!�2�"MF�����X���KV�w<�%2�M_�I��$�OD���B<�����J��`9���)�!���r�¹�P�D*/���2!�ah!���#S_l$�f��dQ�ݒ��߂*L!��F
�L w	�zE���'�@�H�x��#���P�P��Sap��M:L-���J`eEx�O`��'=�)� (仃'یBx��"���6�˰"O�q@�	��@�aKb�1h�Lm�"OaP����`��\���3��"O���lr��-�3|�z)�u"O��vJS�-��H+A��usp	A��>i��)��1j�L�B��ΥjՈ��1��+���'*T��d�'7B�|J~�A��99�p��G�fp�3�C
Q�<Y@��d�f�B;R�&D�S"ML�<�#ۼ|����#��(���H�<)�MםB���5
�=bxD����G�<1�Ç�;i��aڡb`�Ց��^ܓO���u(�O�=�S¤�BHC�e �s�۟�&��)�gy"lG",*Ȼfc�7hs����)���y�Q^�H��0��#�$��y��O��z�1�
��} ���qAϬ�y(RC��U�?A���I2F��Pxb�)�Ql��\�pH�Ĩґ+��F}Ҁ�:�h��=a0�A>�R��g�*� �ȝӟp�	lX����O�N����ql �Y�b@��;D��SvA�zb2��Kߺ�
T��=D� 9`�_�#X=R�H�8����'j8D�8���_���K��X�Y�(�RT�5O�DyR�G:nJ9XC�+����W�L��~2'��O�)�Oj���>i#�\��:�b��Ǒ8���k6`�V�<�fM�iH��&k�T5P�Gi�<y��
i���uA�&/<�� �Qy�<)��8
;�9$N�Y½�eQZ�<�O�3��2&
�ڵ��QP���k���O$�9j`&15ʱp%a�m����I�h��������v�)�i	0�
�ː���3^�M��LGk+!��;m&yBQ͓�`���k��H!�d�,PD
���/�|��Aɂv%!�$
ZO�9eD�J�΍�s
B�!�$PGS.]*��;��xH�jqO��D~2o�:�?)�O	�s�  ��ڙpmr���[��R�|�����I8)a�<�7.G3@O�t[�/�Y�C�P�2��¨-��X�΅=g�B�I�x��u��
�&%^��#�
�T�vB��*H��!(9�`"E�^�hB�ɛ0��!�@��� h�BD�H2�Q�'7�-A���L"<�X�a!���C���&3���I֟P����#��� ���9�h��(�+T�B�I�-m^��qJ\�{戔s�/	�ZB�ɸT]&� �Q��\�Ї��LUXB䉌v�>���Ã6Lh8��l�p�J��D�q�'���c��ƙ��%P!�ۢ��(q�'�0�K��4�����O��[�$%h����$u��	��[�$`���&�A� � Gt�$5.]�t?F�ȓ|�@9�e�-Dy���L$A�bф�b+����`�����lr�ȓp��$0�&��i�w�>�ܴ�O� Dz��4&ɖyy�p����>'˸@
�����	��š�O��$+����m�����.��"��b�L�yRD-k:i�4O�.0E(%l��y��X���놆�
}\yQD'˒�y�g�m}�p䃏�z.*)�����y���==u��AK&q��ih GȊ��'*�#?�E����ܓ�L�hFa��]8��!�=�?AL>)�S���'(���Z#��hi,���f��MG!�	:��ѡp�Ĵ3&|���R*!�$D(7�习���@Jm:�A�Vv!�d��>�p�$ =J��9���+#�𤜠
�\+%�3y��D�G���m?\����
=��>q���^ j�`�v�Z{ج)!���?q��>� �8�G�?��L[�"�)b��""O,����s�����E�<��"O���QfFI�Ѝ��:{*�Z"O|��ä:/pCs��~����'B�<�ޯW5� S���2.�H3L�{?Q��Fe�����'N2]��`d\M�֨H�@�!qg����:D�(�GزV����j�+��E� �#D������;%���s�f�$.A�\I®!D�TK�b�+0���딡!v(I"�>D���hB��(��EƬ8�<�!u� }"�4�S��L�����J�/vJY[3D͜<�q�OiIAI�O���3������8���Y��Y� ��������y��E���[�G��jP��!Ð��y"/��x�P)X�e�H�R!�Q�yJ^��qႨ��a �1бnD,�yBeܜyd�� ��*� ��@�C��'�*#?� �Ꟑ�g�J
�pt�2��4�>l�V��?!H>��S���DX�^�XCB�Q,�$2S�]�,�!��.�B��#$Z:a�*�w���W!�d��~�U
Cd�=H��e���v�!�DM�(������E,<�Vy�Cm�F��ā+M����G^
xL"6%".��$�>����X�s�, �W�W�}��5[����?9���>I��� ��p�j�.c~��R�cGS�<��C<o�y ��w`R�+�J�<.�Qھ�Jć!�b!�*E�<�2 �gm~�`Fĝ`��;#d�\8�H����-�L�ە��> �ݡ�m�F���I����\��Y}��Y�5�آ����9��9{����yH��E(
%Q����4-�Ա��yB���J�`��)�$4RJI	����yB�[�g�X2'm&t�H8�hO;�y2�6Rzp��Ag�@بCoA:��I��HO�$�zwΚ�����$}}�=��>��֑�?y���S��q��yC��1S��Vi��C�	�N�NhT�X9T30��Q�ˣ8�bC�ɆP�ɩ�X�"`n�(�+�%tB�I���B�aҀ`
t��E�I�"B�et@�@#� ����G�U��X���<I�� cNxԙ�	J���:U�C�4���%���O>���M1��%?|8�a4�������E����s�Iy�G5�&m��[�>1�5C�D�Xu�QF�"��ȓJ8���J}R8�3D˺%����~��m�5L[�\��`6���҂�#�#<J8G���
,�(���:F�x��Rɨ�$�O0��:r=��@�շ9��Q{�M�@�!��]1 ���q�+�9`E>컕k�NK!�Ev�iP&�%Բu�a@Gb,!�_�vpi�CV=��1�i�-%��xR1� ��M�pk��<M24⃋��\�X��$�"Fx�OL��'���9L�r�&��v84��H��$�C��$q��
Ѩ�9#fԨ�j@>1C��"h��E��/לA�����%J+�B�	Lb9�ÆȀ	#8t�V"�x��C�	�q�z0�e��#�|5oZ!P��'�"=�z����2cj�Ј7�ʕ�F$�R������OH��-��	V,MQb�ɍ�3�24A��5�y��٤#�4��#w�H�jA�Ҕ�yB%A`�V%�q�Зo*���
��yb*K$���΋�R����m���yr�B���\C��#K��$C5����'�l"?�rʟ�˳��8D~�� E�MF8��O��?	K>��S��򤗗g��AB�˾`{"(��Iս3�!��  1��e@u��8���H���@"OԌ�e�^�2��KE���+����"O�Q2+_�F	f� �H�#�ܤJ�
OV�k�3+��2@@��8��e�����O��H��S+�~ ���ͼHqh��v��!+Fȵ����?	�	<t!�̇�: �A ���E�4��ȓF��dՋİt���Õ���q�����$���7(ܣ�����'�
@����+O�UQ�*�Qo���r܎- � ��I�(OD)Q�*�)>��y�5�Y>}~����O�rb�i>}�I���'\���צ�1�P��-P}R���''�e�T�;n�z��Oչcb���'c����f>w�j	����X3�1�'x�`�􇎋@.��%�8f�t	�''4� �=/z�B�.�3W�>�N�h����)&U
n(z��N<3A��IK����|�����?AL>%?��S�T��bP��N��@���?D�$�f���T�b9ص́�?U4Aa��>D�hơ��b���'#˷Q��v>D�V٘ ��) E�s���	�Z��y��Y��r㨚(g/ tȱH���'��#?�0G�ן��$DٚR+��3�Y�&��D��?�M>��S���=4.� �偙�s�0%�r�X�E�!��<A��#wA�9��h3��be!�S�c�%�%Y�v� ԩؓG-!�d.]T��4�hr�`M$���Ȼ.������-7VP�1�D�_���䑞u��>	sg-��"�u�2��!���7똰�?)����>qV��
&�(l'��#iv�r�jc�<��aA S5Z�颥�\�>��q�_�<�aP� �n@�6��$����K[�<�C�x=\H�&�P��0jN{8����dF�q��)�7G�b*����L�/����n���ϟ(�IC}-'hpZ�
(!�[*C����yBg�0�,A��R8&�H����$�y2�Еf��͛���+"P>%�!�\��y2��:�ɥ��lr�@p�ۥ�y��Y�"�����m�+Ro�� ��3��	?�HO�2��4�S:\�ҁ�&$s�4:1�>�0�ϵ�?i����S��/�ё��~\ޠp��Rw��B䉝2�8d[0΄ifzR��bM�B�	�p��a���)C�j���k�Am�C�2i��5mޡoX�Q�gŏfKdB�	4%�]H&/��IDT( !D�hJ���r���E-/��8{���#vî*T�ç!ͤj1��d>��O>�|��������pL�Vc�=�y�ȓbTȁ��N����q���T�O��#*`88soK�F-|��g�1m�,�ȓ��e.؍\�nMb!B+=L�a�rt�G���;jd�!�V��e:�=��r�D�Td�]�8<	VX+8�*\��j�/XE4���O������t}�DÐ�:z��!���M�!�$D�g�����?q�8;�-g�!�d�U��i[ �F&�ƌ"�m߬b�!��ں�Kg\;� �6Ώz��x��"ʓ{j�P�S��)��a�D�5W���E��Fx�O�B�'��Ɉ8�
B0���!�dJ��g�JC�ɪ�AH��ep���GKǋG�.C�<7<D���>�Ȱ�7!B.Y��B�	�i*���M�Rf����şz��B�	RYРs��P�P�wiɸ ���'�^#=��얶g��m9T�X�	�.��@cQ�D�7� ���O��O�OW�s$��)b�����?&��'G�P�&�"���a��,A���3��� �]ytG[�7���V��To�i�v"O4P�P!M{�h`���h_���F"O6I��*�<6���냁�E^z�`��d]�'�fX"��V���R��T�l�%���Jb�vje�'��'���Y����,J�,�@���ܖ.X����*D�� �mδ��S�Z�65�'D�@c�b�*դ�%��Mʬ*p�#D�|���A�,s�$Zu��k�֙�'�+������v���IcN:9�T��m�3XQ�$�@F0ڧH��Y�)Z�Xl���J�J���'���'�~���$j��`9�c��z�0	�'aRX��e��$��Hi��F-Y��1R�'y�Y���%}�DI U�?_h|P	�'�f�
&��F.�]9T�P�Z6�9�
�Q�Q�{��s�u���"i2re&�i�'m�Y��h���O��V\�ؐ���%R�t�>o^c4c�-~(�k��OpTR��j�g≽[т�H��F�w�� ��@��Y�v+�6.�`j�'R&�A��4�3�$�_ Y�%F8�$)Zi\�|��	y~�jҸ�?ͧ�HOL0D*�a���8bH��Ft�4"O��vH��29�g&�\2����>���i>���_}b��h`�hrV@O �zH�m^�I���
������䟀'��O�\�("mV�{�DՒ��ז2��r�N����4OP�{[��X��'�d-P��ҽWh�a��s�h��Eʟa��]��8�J$�'��	��i��?ҙz&��
L�2�m���?	��hO�c��(6�l<�|��a[9��Bi9D��4 X;��sE\���Q��`9�	��M����'k�����-`d��BW��Dӧ�V4=���'1�'��Y��!�{Q@�Y�'�<l{BJ:D�h����355�����	WB([% ,D�(B���i*lAT����iiG�/D�������L�Y��T�&3ȕ���.�� rFD=�<���`��C��1���LdQ�(��#<ڧ%�M ���]�Dmz� ���1)A�'o��'�ڕ�P�H
�x4�n�@Й
�'P���j.X�F�B
�{�@���'�b�Z�m�O��m;�I��/����'�����t���� 8�(�Ǔ_Q�D ��!\<��d�m`���Sͮ���)��|����?y�O ���h�-eڴ����L�1&"O0��Ӥ� {v�q��øq)e(�"O� �2͛1���րQ�(�4x�"O@����$GM�[��[/u�|��"Ox��e߭lh�QP.G��p("U�>QT�)�S ��M�*�h�´���=����wb/}r���z��'ɧ�'>/�J� �7=~th�O*�,��zLi��L�j�x`�u�P3�D�ȓ�0��1eӘiA���g�?�\��_��*���K�����+r>1��M�BuҦ�"R<f��clм"6܍�=���I����$�<C�!�JE}��J��"VzBL�Id�I�"|�'���vDL@�pPq���Z���K�'|X�顬�.JM�)���E�R-����'��H�B�	 P*�B�K	�BY4��	�'FŃp��3L��m�$�B�:��
�'\@@��ӻ+6�Q	A�ۡI�0�q�{�'W��9�'_�2�����7$zj�)�K>pQ ��5�'��'ߠ��2*(���lY!zc�0
�'�\k�ǖ�pL:L����wt2MB	�'R�7�Ļ5iʠ �l��}8@��'��X�_9�T�ʡ�F�!���ǓQ� ���V�����(D'�p|Ȣ�3D�����  �   .    ލp�F˸��%�R(O5f��p"O��Q   �O4���k���W�ID�4��B��0<�bH�Q���   ;    މ04���R0�Q(O5f��p��'l��_��p>���   ����XѮ1�'T�����   �   ލp�F˸�41C�:�1�#l���_�)��ToڬrN�'|i�@sļ�M+�'�����Ď_r�r�K��<��'؛�c�����	/
j����ο��rӭ߳G�L	�@9]��#<ɶ�k��4��=(����&$�4�ӳ��]y2L��(����DX89>�ݺ�4=���K���N�z�^@�S(��ܖ��<1��V��O���6q�l��'�(��S+�D���x9�l��'<�]kfE�a���	"�4y5����'.tL@1h�h�r��C�1zB<��'��*�N�+A˒��p����'��H�k@�@c�,CD�`�P��'w�=�GWTI`[QHD��4�J�'�:�pK98�S�/ո2`��'�b ��I�}N�u��$��q�H�1�'�I@�"�%<�1��\%q��c�'/�LK�q�(�k��Tp5�Г�'p�����(��1i6dعa첝�����	 ����$CG��q�O"���'}�Of���>�F�ѦI��~��0��.C�m�$�q�&y�=q�+2�n��'�����U�����EkQ9�|Q��Od����,�Or�K�k�O*��u��zl2Qg"O�(��  �n-��ðiO:��f�'JX�J��dт8#d�p�S�
�b�M��M�ax򠋄�?I�yrLV�7�|U`�!�9�� ��.�y�V9*8=0�#	,3� �H�����?�2�'PL1 b������h�N�MX���ҫl�����AC���j

G:Ÿ��[6R�u�������	0a��$ڣϒ/*0,lBE�¾l.�B�ITQVm)�D�w��ѐ&�~NC��-+�����(��[��s�+˿0K�C�I	\̀�'�.Y�XMH#$M�?��?��퓨)c�A� �Z�P���O�!!��ċqO��S�� ��z~�i�"�V�9b�A�]��L{����yBI�*.D�� #S��+�^�y"�� �k�ፇ6:���y��M	���D�%/��0�R��y2�Eyֲ��Ќ�25�p�%����L��(��)cL�*b�*E���"H`�3V�TsDK���\�)�3&.�p�_��PU�HݮB�Ɂ2�����e�*Y�@����O��C��sy�T棔(H���q�ːl.FC�IZީ1�f�,�[��ȯ(0C䉺I�
Ĩ��H? ̑�%J$!���O2lE~��M��~B   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��R&�4*�ب��P�R�B��eN�uR/�P���N�G(@��������� �5   �  �  �  �  6%   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�U曞@�VM�P������@��P_`���'4r�'d�|J?��f�s^hy�&A�x������ b�8�`XTv�|2���,�
�*��ڹz7"a��iRȖ:[�Fi��	�[ڀ3�F�\l����S�
��0ɂ��O��d�O:�d�<�����'�
�y�H�<_�^|��'�*�$���'�j��ULT1H$�au�C�'O��k�{�eӼ���<��E��?Ѫ� yY�"�9K*��1���+D���ϟ�'����?y�a��o�'��T��ȍ0D��,s6a�D�0�	�@��i8�*,���m`���r�ښM�媓E�w(ay���5�?9�����G84��������z&U��oÝ|'���O`��8�)�Ӟ!KP����X�t��xP]�K1fB�	/Z�x$KW��yL�X��X6y{�� ��(�'�(P*4�c�lXPO�O֓���]RT��1�`���XHX݈��'�K�8�2Q�p��o�,O��;��ݝ76�T	��44։��xr.G.H�(*�* LgRd�Aʎ�F�&?)`q̔~���QA�D�>Ģ3�2�� 	�'��O��O�Hx��D�D����q+f�pL�D�'4ɧ�Y�rql_c1Z�s$Lu}J�P�/O�Ilǟ���ß��}� YԊ�3?�,4AE!KZv���'�R�8���O���O��Ļ>9P�˸x/6]{�N���j��OX�9�|��ɑJyj]�Pio����a��n�c�\��',,O����ѕ4�x�
��)	��i�V�Oc̓
��y�)�3��
;v��#-�]�K�K�� }!�Dʕ3xȓ�1*L~\ �O�e�����E≴Lx�Hk� ��g�,� Ŝ�mH#D�0F��'pR�'��I���I�|��KӬ2E~M��/\�d�L��MB6���P����>�@ŧ�fD1+
A�p9�1��㊴K�.����>Y�N��r� �O2e��
��,פ���؟����Ж's2��êv�K�ƒ�\���Z-`�!�G}�pk���	&�Q ��BiqO��nZ����'\UZ�Nw��4�i�>l"e	*�9�TDC�"�t5�a�C����'=�'e�� !r|Ε�2E&}��7s�R�/A����g����<Q'NҞv&ZJ��
AJ>L�Fz��èVU��I�',Od� ��'���' �HC�	�.���o�p �C�Ċ�<��?���$�ߚR���eNC�yq���'B��Px�R�,1b��)�[����5JC�Z�����'��O�9����Ԡ#ň� n�0��m�(k�B���DM�����TX��T�R���0-L�G�d	�W�&D�����ʜC�^�i'D��7���+��6D��`�$o����S�-������3D���De�w����-�$[�D=Sv�>O�!FyN�3T(���V���Y��ȓ��ύ�~2kB�O��OF���>� Z\1 �Ķ,P�i�	�a&jIk�"O���ѯ`��R��G'@i"O�5�D��6s�Uy���p&�-�r"O�HGF�>*
���DT�:o0M�t"OX� �l��E�H*1��{�>�f�)��t��,�Ղżj>�Ѣ�V��Z�'*��ҵ�'y��|J~*�j�a��u11I(90��B#��o�<Q�ey�� h���"k�Ԙ�hOG�<��W8�,�宄�XA���PC�<��E�+X:��څm���X�e�C�<�f���� �]�k����~�J�����G �OF��b�V�J����FB �Ԁ�hDП$'���)�gy��Ħ-L�|0��[1M(Ȱ�֝�yR.�M�`���Kǃ!oP���J(�yb�)][2T���cReO.�y�hއZ�zD3��Fkhm�b���Px� \�@.��Sd�C?Z) e`ݛfѶ�E}����h�P��ħ9��a���^;z������	BX��[��K]0�x��]i�RT��k*D�0�&D�uN�)Cs�d�á�Զ4R!�$y
�)3��n����W!�%C!�]+�x�A���p=�dm]5h��xR�"ʓ
>�(���@P*��Ƌ��UT��{�}Ex�O~��'�I�C�p����D�np�-�DيӁ;D��@��C$x��S��q�feƦ-D�$I� ��mq�]H�)O"8�b��Ӎ9D��i�S����TY��3D���4)��K����у��kY� d-}RL8�S��4F����ɆS��ɔ%�74j�h�O ��e�O��*����'��*���E�T��a�*̢�y��F�iz|d`rM��S��l���΋�yb�k�(�R��/ENT�)B@ƾ�y�G
�bvXHi���&8���*�b�<�y���o]�,�W`�&)o�AbQ���'?�"?yS�P��ʧď�`����(�)K�8����?�N>�S���DW.'׺�&�1KB�e@GZ�!�$X.���q�I� \b�r��mt!���3Q�`X�bQ�q<�88���k�!��ֽR&.)H�A���F+V�~(<A���
x;��y�	B�6Y��m�-<�B�>y@,�b�O�*�2�ЀZ-T`�J���&�t��O���#�OD�a옳
�d���,�� ��H�"O�Pa"�A�>��1�˅����"Ov�����!�P!2�.Z<"#"O�i�l��9=�(�ċY�:E�+R�'��<i�Шfqm"��'
L���s��k?q�o���4�',r_�|�¼h��ZBh�0,�޵8��&D��r��U��u�$狡7�53�b#D�\��
̦T
|X��NV� g�\��K D����(��`�̆�\��dK2�1D�`��nA�E>�0`5 �D�����/}2�?�S��o�8h�"�_R�T$̎C(E�O�Y!���O���?���( "���p�L�b�������y��@��q��۳_����e�(�y���h|��9��;\$�T*�H6�y�$F6_�V�yCm�2Y!�C�n��y�\_��*�SP��'��"?�c+�ן���57�t�v`RnY�d�!�?�K>�S���D�^ʁbъN�ur��P
�H�!�$��P�L��	�:A�U"_�(�!�$��:����P��VJ��P�!�D��e�f@�3BJ4&P�3�	�j���}ܾ�k1aEQ4�Q��*Q�xI���i��>�#�$��.^d�Ђ昷w�*a����?����>� ��)7ʗ(��A���Y)d�X�q"Of�9$X.%����M������.D�P�@Ȑ�*�q�E�-c�!ba�2D��Y#M� ����T�� ���"O�aDyҮ�2	vq�f�#��(�d���~BlW��O�I�O �d�>���2dK�Pi�j���s�*�U�<y3F *�*<T�́�B�kg��R�<�a��Vf|	a۾x:^4��N�<�Bg�4Z�2��0
�9��@zP�B�<)DIS��V�U�:]rN�;���z�D�Z���O��͂�	 �p~\u�ooW�i�K�Dí����I|�)�	Ԑrb�A��l$¨�⢎L�t�!򤒇H��Xrd�U�>�2���b�<�!��קJWZ�� L��%�$A��Hޖ[!�DL3�l�1�푫H��
f$j!��Z7'��L���S�@�F�HS:}cqO�YF~R� ��?ɓ/=}�����FejlH��ۏ<���|�����I<ˮ�8�b�$��&�@U6B��a��9ABM�6~(���D�L�B�:�x�'�h((ШD�,Y�B�	�W���U�A>}J��k�2,#�B�	�x�����Q=0	"0��f@�:� ���IN��}����T���Tz���F�k���']a}��Y�d��T(GF[/��x6,�?�y2��i��|��ɰ&��U�� ���yR۔=e�:��S��h`�#
�yr�W 
�V؊Q��M�lxB5�6�p<���I-JR�0�^�h����R(C4^�I
�#<�'�?����D�_�@��e�
>�P
�ȁ�V!��"Q��h�b;G�BÖ(�7�!�ȔY�F0�`Am�H!� 'Y5 �!�M�vs�q���Y�\�b��*�!�d�"�BEj*�!>2��'Ő��<����?�!"ܺ8�n���B����]�7�3}�Z�p��'*ɧ�'(3�t����8|�-p�d�!2���W��͓�2���(�Q@<�ȓ�-��q ��Q&l9�q��Q���y�h"Xsc����,�ȓB1��Q�X+	���2ҤX�)�40�=���	�r���dRw�,X�3Ņ���Ig�B1
&��a�	֟"|�'�Й�bm�-N����uA� `5Ҙ;�'�䐒n�g��\9E�,EQN��'N�]ɗ�ڱE�����]f62���'dȌ�g�R�j�NQp��=nH�a��'�8ԃǉ�hf�<q�lZ�P�|�JI^�'c��z��)D�$��t���x���a]pTa�%ɟ��	]X��,]�T�0��QK��pS�S�FW!��=mpD|��ŉ�K�H���,!�DC\��óh�9(�<*��W"g!��yl���Y>'0�����g�xRI8ʓi�����+cl��IE����3���Gx�Ob��'��	Y���c�WsS2$(�dA�aP�C䉧q F5���j� �!E���W.�B��W���i!�H
���ĢQ�[b!��ˑ8�����Ѵ
ڈ�*𫟣�!�ߠ1 �B�e�C�f�г�Q*��_x���?����$c�X�ƍ+TL(�A�2}�!R�(���'�ɧ�'8�2��AJ�.��T�A�ȥ[_q��F�B�@ң�mH�����4�y�"O�yq����,��l���ze"O]���9�E{�-H  �ؤ�g"OV�z���W��,���3K�LM���$FZ�'�B���`�νC�ņ��6��H�'Vڔ��'J�'W��Y�����ZR����R>W�4I��5D�� 6 ��SDݶz��?�B��"O�$
�a̐[Lp="Bo�G3tl�e"OR���C
�b4���0oW�3N@��
O�qaJ%,���A��K�]�lA�Q�ΣѨOX�9��S�?�x��_ ��L�di��%�(����?�	�<`H���]��� +"�\��ȓ)�	�v�ͳ����%Ʈ^<�ȓW����k�
V��8&�%t.֐��p��=�Č �gԠ�3�,�"�����Ɍ�(Op(T��`�Ր3N��ki��:��O@����i>�������'�.�{�
 (F|�0�h�w�X�'"nH�$Yu�xEpU�D�sLZt��':���jZ�a&4᪄J��4�� �'����iĹz:~���  ,�@�'~y�G�^�#Hv���@4n�~�KL�ٍ������ 4:��Ϊ	I��Hy�*�l����?�N>%?#�G��L��<�� Y={��2 D�x�$풋M���X`f؞hd�}+��9D��7�D5�P��p�"|�xQ!;D�$�f�\�J;�$�@�۶g~�f�8D�`j��Ts�4E��F;�ek�L*�I"��O��hu�'�RQ�!�T*e���(�4&t��Q(�Oh�Ov��<q��[U�h�� ��U�\� ��u�<1E��}~z��1�dC<�x���s�<ip�?2m��XPnL�Jd�@[!��5�*|�&�H";�	b��5o��d%Y��s���HƤ(0e�55�\�����8�>�1r��8<�p,�d�S	_\�B�I��?�����>I%�9�(�`@�U�;�*9��o�N�<	��ю5��9��*[�vIO�t�<I�Ǌ�2a��+Ёds��Z�+\�<!��\�iF��MI�}߬���b8�X��jP����;Lq6�?h�dղs��������Y}�.׹Z��ir�ڨb�n���"�y�.�$�����Xq�8���8�y��ۛ��#`���p'�Ы�y�eƐ�Ψ���Z�vB��qw�ފ�y�)�yh���Z!d��%��'����
�HO��X�G�Yv���C�k"�qӟ>!�X��?Q���S��7�*���6^�h���|7"B�I9]f~t�
���5/� \4B�	_�x�"�*F�4�P�f�3��C�	�'2�pa�Ϝ(2ٺ�r��3B��C�Zk(1�� %`��`)��� YE��蒏���.����oT�a�8�tEN�r
L�D7�d�O>�X
�m��!��)m�0 �(�$:�A��#P��c��X�[��٤SNX��a�p]�Q
e��LJ��Ҫ�$��:���	��I�
��4��%v�`�����*K�Ġ��&��|��8Ё@0�%�.\E�4+p��d��\v�$�SBO2#��d�O���Ě*L��)O� ���YFF�>\!��ѵX�-PU��t��)b��YD�!�DH��Pl�CL��x�.
Y�!�DHs2us�ԾS�*  ��P�x"":ʓ ��Q�P�ܮF��,��
�,,�(A���Ex�O���'�����R�%o��ܸ�L�?�B䉑&h���W�kr�tbE��<0H4C��(>�3G�F�W6�4Ó��AFPB�	Z�&����jA'�$B"�����!T��r�̈́�G�0�
�/-jx��>��)���K�8Y)��)D���9�`�7{�2�'w� d�'�r�|J~�";jS~5xS��->h��Em�w�<�7C�56DD�� *��Q�� �av�<� N��da��n��([U�I�K�B`�"O���"A5S�t�jGD�Bt���"O
e;��_Bb�A�#��
V6�ç�$�z�'����V�H�ꄯH�N�8����%���?�M>��S���đ�c�FH
Q�4E�DT3��=M�!�D��7a4��!��[U�(P���!���� b-�v��V ��\�!�d�"�i ��]� �ZwI�<Bɡ��N7�8��p��A
Em� J�.A���d�o��>E*�ё2Wz�s�Qh�A�vhC$�?)���>m��+m�m���Q�F�$e˂,�F�<i�(+�&�q�'�nڎd�C�C�<!R$Y03����  �'F�w�<�$��U3�a������h�v8�0ۍ��p��$���6%��rjJ�pB��-��UBZ�O�2�'���+n<U���� ���2E��
sMC�:]C�kϋ�?!6�'����'5Ї
��?9$ɀt����G��m�
� %�ȟL1�������oZt����,O,leZ�߈"h�t��'�	>E��4�V"=At ��Э[�	�$1r�a7��W�<���ǟDY����,�
�Q�WL���{�����'v�I�vQl<iR�2	�8 u �ycpE��\~�'�2�|J?AI2œ;EU�u���D�8��jN9N'�"Wg�=��� gJ�dx�D[�)(R�T���\�R�جb)�D�`L�!��*��K6L cx�P��ʔ�mz����⃾ht:�Z`�C�o����O\�=i�}�cK�k�P���kWJ�,h���إ�y�c�4~��䃖>f������'�6-�O6�	����i�5��i>y2�'=:ހ����p?��b�c�Or��?�����t��6����ݺ�D�OA��PBAԖ&�2%b�'��%l�j�.r�+ �3 �H6��+3p��݁I��Hr�+>���J��T�?Y���$̇I�VH��Ћv!Z�pFJE�h�qOh��),O������b��U�q��Q)D
OvW�>s�Y��L��?o @����x˒�;���' �H���w"J+�M�5��:����.c�й!��O��8�OHesv��S�Tu)O�=xJ�,��"OF�c��W���!�X!"�HQS"O*P�ǉ�MLD�xs���W��`y "O�t�Q�J2n~�����hi��j�'6F�<ِ$F<��(7HP�@g��5��o?�@�G���$�'2U���v�R-ip,�G f,��@��;D�pC )Kn�V��t�:�A�2�4D�{& A6 �J��Ǌ��m�h� D!1D����V5n����BT`�0��<D��yVR$&D���F"��g�vܩ�<}2b;�S�']r�0�#P�3�\1.��pF�X�OV�C��OL��)����C��ey����a���[u
��y��D(Kk� �& �&K8�(���ҝ�y�`�v��m��Q�ɃЄ89�'�l}�� �R�x�a�y���
�'4��i"-��G(^��`�Q x'2�ȉ{2�/�3ǌ-�	����p�"yTh�c���20�����?E�,O�)��cF�e<JU�%�/!��1�s"O~̘�B������] |X�t�%"O"͓F� <�� �lH����"O>��U��0w-�D�����YL�12
O �G7W�ى�.9{��=�ꐕϨO�����V�0�tO�5;����qO��j�4]i���?1�b2\Zg���ێ����Z�@�ȓT�pd�tG
�W�p%��8������%��`K�R��b�� 7S�M�ȓn�bUs�*ްT�P���a�aLXQ��I�(O�ɲBOC6 ���9V��V$��`"Ob��A@  �@?�y")��~��]�?���V����y�+��R�b���A�=A�Ԋ����yr��w����&�K�t.�+�y�oH�,��R钀v�"%����y��to~��%��gθ(CmN��y��N�5��9P����i�Eϝ�y��_)��-yŋ��J��Ò��y�A�4L�#�ܝ�� ��y�F|�u� ��t�T0R,ۊ�y'� ���)n�%r�9q톦�y2 �:6�up�/lc HBa&�$�y2)�.Vv@�F��-~�Z����y�B�(~�xCT��xy����#8�yB�=�"m�w�*_՜ȋa� �y2�Y�gO�\Y�j�Y�J�@H���ya�>{ؽ���'�A)0��y��7�j�q�kO�J?�`t�
��y�B���@ D��:20ś mM��y��!����f��+:`�I�gG�y�&��,�bE�w��05t�;�]��yR(U*�D�eO:u�1��#�y�k�3(������'J9:���y�E!ɪ�`U{���CO��y�!���̚��	t�|@��M��y"-ϻ"����b��X�>�顈���y�OW�^���P�o�:GR�Hi4F��yB���>�ʤ��,�4B�h��"��yB���� xF%6�B	�Ʀ���y
� ���v�Ę�B$�ԥ)�f�@�"OVi8 ��6pR�K�>2���i"O�I���F�,�l8�c�:|�p@R"O�8� i�.x��i�X�b�
�"O���2W���W�M�(@X�P"O6	z�
9\��ZP��$K:�}
�"O�m"��Ȼe���"�)d{�Ԃ�"OjWnڞ �#0�ҵudvHs�"O��A��֘;
ȡO�zD0Q��"O����!W�\;�MS!D2���"Op�l0"���1��O M�~ �"O� ��2H9���89�ԐSf"O��)b�W��0X�Bk�7,�
�s�"O|P3����������O�R���"Oru��*�zP�<�
�&tEJ5�"OPd1�N�w�J�ǋD���u"OP0�D6E��!Rċ!i�f"O<��'�ر{�Ђڰ
�mK5"O\L�B�J�sp��VK��t�hm"O�� ��!{z��SJ[�v1�	b3"O.��SJٰ䥸�nĂ(:�"O��ࣦ(H�V<x��V�xU"Oj 0��λkچ�ɦl�6;� 4�"O氉 �Al����4kN�S_�a"O�M�V�Ҟs��T��W8YAK "O$L�o҂x�6��〙I�1ڄ"O��ѕHh��0���ķh�N5��"O�U��a�"D����ˉ$_��P�"O�`�	ܴ=�ʳ�L#\��]�3"OT��F�+�)��l�*�"O��6+Kw���0�٬�x���"O>��q�.�p�+5��?�~ݛv"O`q�`W<<�l���>`�ZX:�"O`a(��=y����D#&����"O8|�ׯ� I���ڠ�V�?���8�"O�T�P_��"���0k���v"O����[L���1f��a�"O����+��M��895�y6Ʃ`�"O�J4h��n��AP�c�`'�Q"O�q
��֯Rv�|�g���"O���� ۳v�,,{�Y�R�8�"O�Ö�����8T$*����"O�\�d��L��l1�d�>Vh�]k7"O��@K�<k��a$D�-EVD��"Oؠ; �?��,Ţ��+D�j "O���F��X}4�H��<v%��c0"OLl�ueS9F���RkA�D0�;�"O��aF���LU�L���<^��p"O��0��W�?$4���+Ѣ=�BP��"O�D�s/9$Z���%��q�ݛ0"O2H[�b? �j�;�&�Lmh#�"O��"g�Lˆ #�CO.\N�;F"O��)�d�*J�tAT�ZgF���"OJ�I��C�6�Pxه��}8
��g"OTZP��)h&��o̱)�4ằ"OuX��/Ww��(� ��>�P�Ib"Ox����,.pP`�� Ա"O�-�G��+��"��[�ԕhW"O�\�����~�8=J�J�(0�Tѣ"O��K%��z�zD���N(���"O�L�p�)!0VA�Dh��-4"Ox=�Q�N����RG?ZK�Ч"O�qhVI\�R*J�buE��$Ap�ڡ"O(A�`������S��`�`"O� �Y{&aO�F��(��ԩF���A'"O`��TD�1qfxY{'��Z�1�%"O�T�e9J�vi�g5<��=��"O��"A���S`d�bd`�XWB�#%"O`Q�N�I+���hF�1��峓"O�Xx�+��q�@<��GZ�J�,�"O����-�J�65��� "|x4(�"O�< M	;9�̙��Q j:0�2"O��p ��\�����)/��@�"OFij��� %|!���X"�Db"O� ��J�^)JP�e��+�h@%"O>�4�SP�ᚷ���I�p%S�"O�q�WDQ9K�p�DeQ29 ���R"O �jDB�-ɳ���7����f"O��+�2�0	��V$	��0��"Ox|ZҤ�R��"�a�#�l�۰"O~�Ј��@Hk���7�D���"Oȵ��܇o� q��/�_���I�"O&��D���!�|AC�8��u�"O��p�ѫ.~��2�N�%{v�;�"O:�3 �)!𨫲��0z]�"Ot5SHF'jޠA�D�l�ж"O0 g�m�n�0T"�8r��ur"O�Q����V�Y�$k�:a�tL�"O�iS�ڈ&� hr2�H�V�B��p"Of$�LP�"�v}dL�
{���"O�&n��e��(�G�Y�	µ"O�D����;|Nq��&��Sq"OҘВB��/��u��F�<|y�"O`��s���/·>��7"O4D���5J�x�0�`��_���v"O�c��� ��S m�}�@Q��"O�����QHhJ�#�e�.�� c"Ob�CeA�!�2��F��F�: ��"O&�)�"�r\0�[�d���Щ�"O�p�3��?<d,��D
!F��x�"O��N�,��lp��R%s!�\p�"Of�:Q ˙;-Z�7�_%�cb"O:܂S�ɷ]�w ^�$D�X!"O�,�C	��>�� �IL��P��"OD���L�Q&��0F� S$"O��ӄF(&�uȦ�����z`"O��q�'fU�#����� �"O~��g�\���ӂ7��;�"O4��¹��)r�! }h��G"O�I���G�r���h^��"O��)H��5c7/�S&�A��"OV���A!*\��6�MzyP��p"O�E�s�Ϊ3͜�*��ݕsr�y��"O������0$���R�=({.�P"O�`�q�֝u�Y�2G��Dz�(�"O�����u��"aM�w��}��"O|���m+1���)uZ��ei"O<D��aϋ�a���G�Xq�G"O���k�N22ǈ��+�"Ot��3ʐ2&�䐣���"`����t"O6�xѭ�0K�.IS�/E�)�hp"����zt��͛N5YvM�^i�'�����[l��E�B�N)�'��g�*ZV^���\&|�X`8�'�ܝ�ơ/t
=�c�߮!����'��`�3�e@L��"n�i�X�'B���t��=W���#aoG�
G��	�'��M!�"ПLN��0�>L`����'�����	o_�{�.ԏE���p	��� �T�4搥!��Q��='z!�P"OR������kH����>3|f�pR"O�]���S�.�>���"Άdl w"OBx+���U��dK�2PT#"O`)B���UM<u��ȓ�1J��ɕ"O `�/��y`����|��"OL�������bv
�m�dt �"O�M�A���"�pJ�&	���"O��SEFN'�Ը��c�a�:�P�"O(�2e/՝
�,�r�kP��b$"O�4�S"Ӂgd�ٙ���unt�"O�u���E=Y��o1p�-�"OjPX�h�-\��]��i�@O -�'"O~���*E�W�di��/X�6D�a1&"O��h5�ؐ?�zՎ��\�r�� "Oq0���"p<� �������Id"O��+0,��i.��Z"E ���@R0"O,����!7�\<��AB�u���""O��(�KÙ[�fQ�R.\33���"O~�z4�?S���c�+�$lj8�U"OV1�à��x\!%�#1��A�"O6��_&s#B�u��6�"OZUJ�`J��tAk�F@�Mp]��'sj,��b�,Xb�yjg,ߖt^�Y��'��X�����Z���
�LB�~;r� �'���a�lҨSq^��q$ÈHiLPa�'�)Z�hP����4���.!@��'�����њhQP�2����'�t�)D�Hj�%�s��7*c.l)�'.TtS!̢ɺ J%
\q�'A��s��A%B�ATj�.��a:�'̩C��t���┫�� ]�,�	�'`��ǂæ5�����W�.P4�I�'��Lծ�;�9!I�)[(@�'���!���FgB�|�j�'f��+/̥VjX3�#�9�P���'�<��C�_�x���gĴB�L�'�8�@T/:�D���.�K�Py�'4Π# BѠ��Q�C��-0=��'&��1����oI�%�Ȑv]��'za�	�ZfB�����|��'���B�"DL�9ϗ�M.$;�'w���Ứy��С挒q��r�'�ZMyƃ�O���a`XY��T�
�'
�	�q�Q6�bq@�Z�[:���'A�e���<����3���pX��'���F�D����2(�*=-h��'����" R'N���B�7�l��'���CM�8���+A*�%
�'5��AC �/\uh�#Wo����'G���N�>jװ�4��k���S�'�\� �ZC��-�h����'�b]ص��z��k��ϓc�f��'��)!�dG25�=R���4\Z�'����RH�4l'($A��S�"��:�'�`�A�'ϻ}(��4!��LBI1	�'i�*�W.;�:%#�G
.H�r��'��a���	!d�Pr Ʉ�ډ��'��u��&�)a���ʆC�kf���'l���G	[�=���ڑk�2�n(��'N:�y�	"���B%s'&�k�'��	�2م	�P��p�^��X
�'&pyO� �"]�!��H�����'T~<�Ύ�/{"-t�U{��(���� tlu�L3q{b�#Q�@b�2"O���Ưv}4YB�k��
M�)�"O�� ��	4�>�EhM�y@�m[�'XV4XtE�2c�;�EC�_�fIy�'�� �鍲K+\�@�]�
<��'*I#�T���V(2M�2)�
�'Z�b �?�8f�V�Kj\j
�'�:mH&�M�xy���߼RP�u��'B���W��j1lLm�E�'QșQ皈R�vY 1d��.��ap�'~&i��,��ԑSuF��-��J�'���!]);��Q�']

�	�'}Ԑ�����@�`�aԋP�a����'ȡ��N��%�GmZ'`����'yؼk@H
�1�`-Br��8�{	�'E�ٸ���"�M[%��.ZJ��	�'�"`�Q�[	j+�� ���"AH�!�	�'� �HB�)<y�@�W�7A�Dlj
�'�jq�kY9$�(���̗v�$�' l�rO�&-|����A�;h��s�'�Aȷ��7utB�!!�ܞ,�$�@�'���C��^�~�H�bJ�$SF���'���i��_Z��� ��*/�v]+�'~����A6� h{ B�p��)��'ڪ��]6�"�X�ϋ3@��'��[P�T�s�	sǊ]�4t{�'2H1s��A��qҫ�*Sg��	�'Iܩ��_N�xy�'@HE���
�'ۜ�;d�y�\49 B�0}��
�'�9� f[i��M0e_;dxP,3	�'2����	F�8��B,U��|	�'42 ��TÚ�SE�Ɣ
d� �'w�P'%Ƀs��|�g��9�eB�'�
��
�I3@<�I-��a��'��Œ�JQ��`C�1[�L�[�'�xa�5��t�D���^?%G��y
�'��b5K\�5������#l�$��'{��9��'�z�+ �Ȅ:5�e9�'�����h	I!~9p#$�03�%��'��\�����}۲ˇC�_���'�܍��h�{場�WLėPǶq��'#:l��u*oޫ2�XE�	�'T����o׌$��'R�*���X	�'ǆ�Y�KȳXdlU(�`ɺ%�����'���0&b<h��ㄜ�"�ݛ�'x������?d�R��e�H�@���']��bǁ��E���Zb�����	�'��2���z�0�T�P�W�Ż	�'HT�A���*WH�t��R�I�~���' ̬���K1LĞIITf��}M4���'s<�rk��a��Y�ǥ�@�4A�'�@P�N_+F��F�7A����'|XA�\%9�|�Q�ͳu{z���'5<H"�	C�!I2� oSԬ8�'�H��擆-8ƴ{�΀�l��%��'������م���nD�`�~�:�'�u��'�E��mRR���l�'Ih,�Rj��S�)��D9}G��'k�īSl�(b:�)���:�8)��'��4��Ԁ#8�1�b��N��1�'��K�84 �E`�$ۮN����"Ol�q�čGv0��ʆ� � Qc$"Of�!H���	p�䅟Y�
�!0"Or}�7!�Hg�c���2��}A�"O� b�[P�
8x���ʡ!�+X�^� &"O�%�!���xl�S+˶D3��5"O��$�3f�䪰��Q$:�p�"On-b�L�"�*P����q6H\P�"O���e!��az@�Ŏ/"�H�F"O��Q�E�8���2��ز9��"O���F� /%C����ސO��zf"O2�J�.@��J�1�Q�l�B�"O4� ǋ3Y׺����Q#t���"O���Qʎ�(��� '��~~�8D"O��:3 X�%˸��P₄u4���"O�pR�Ɠ(p�����>6i���"O(��`��&a�J�St�Ҙ#�Nxx$"O��b�G�	Y��Y#I
4�V�Q"OFi��/$m�#Q�&�B�z�"O8�80i5G������Z���"OJ���'Y�5vRp�2��;w�x��"O�e�w��s4ʩh���7j`�y�"Odh���O�XheC%��f�Rq"O���N�V��ʂ"C�J8�8�"O��0J¦H���T) ��(;c"Od����[?&��Dt�-,�����"O��YSG�3�@ڕ��!8Q^�r�"OR\�"j�!Ǻ	F�Y�p�pm�d"Ol�CF��>�ĉ�a��4^nB2"OV�@��A=Uq�iu'K)x��d"O^�h�2��hs�fL4_A���"O���4�V�Sp�T�EE�pm��"O޵�W�H�>���ۀA�]���"O�`XfG�=�
�Co_�Y��(1�"O~��U��6_  �,��~V�"O��s!��'��<Yc�M�Q �"O؈(M�=��Pea�<+�!��"ObH@u��$V�xѩ��&uDp��"OT�B��	N�|��N�O~�	�"O��外�S�֙6�SPK�Ѓ"O4�x��;y�&�B�d��5���"Or
��"^�H,��E�.~��`�"O~�5��6d�Ѐ��[�ʥk"O�d�Qa��S��yP��'���Q�"O(��Ė!!!Rͻ�A�s�:�r@"O�p�@J�l�*Y��/�
����"O�q�����A��&&��e��"O��7M�,�p���E�p�D0��"O,�%&
�4�Xd� �U�.�&�j1"O�E�Ŭ��S��� G_E�~�YR"O��Q.�%�n�8"�Q�o�Ƽ��"O� �eڇr�~���� =��C�"O����ޫ'����"O:v:&�Q�"O���UH��WB��tD�)H$�4�"O��H�W�@��K�/D�=p5"O�����L 2aI
��<�|m��"O��y@��s��!`�(e���3�"O>(2H�)��L��B4O�Ҭh�"OҌ���B�PI9!,=Hoef"O�0W䛀H�F�Pp@�ZZ���3"O�m;���+[�B�s�kU�T����"O"�� ��ԘZ�*��L�ٗ"OtɁ�mM�rM(%* ol,Ȉ�"O �������@Fׯ	���;%"Ox(�0���"�4];@���;��������o�l���G�!�4x���"��'�LmS�դ�05BA+I��ح�
�'�j����W�Z���BG����'��x)�"��;'P�1���?'�h��� �jŹlΰ��!�I;@W��v"O�m�d̙!<NAp��:Fv)��"ONp��.�!7���9E!ج�0�e"Opp����r���4��s"��P�"O����i��\!���TH�+r�]k�"O��	B�*ph!G�}�u�"O⩛���w��8��]	�ĸ"O��[�BX��Ph�$�m�0��3"Ot�V�C�(P]�Bc�c���1r"O�����[���Q"��dxڈ"d"O�$sыIg��`��=
d��B�"O\Q$��2D� i ��.pZ�R�"O^U�"K�u��P�� BX�`"OZ��wR�6�Ƀ'#B&AZf"O^�ك�b�b@�#!
�'+0��"Oʌ�b��8�$��> ���"O�]�@�#/(P0�:8�0Q�R"O������*��|���X�9:�"O���/�� �V�1C"O4�)��n�[�`EmS��xQ"O�:� ��j�<<���#�嚅"O%Ň�89EM\�r���@�"Oq�bZ./[�HA��R�XA��"O��yH'W�|2F�^,�Yڶ"O$A��/3��4�7㑦j��""O�Ջ�N,l��G��u0i�U"O��҂�6NX�gAC-M$<�!"O�u+#Q8$��p�Q*ZN���"O��)��ň�!�GW �iS"O&�jvf�'EXx��L�s$T5��"O�X�!��е����;x)�A3�"O@���'hE�t:��7J#�IH�"Ot���N�IQD��$��m
�$�1"O*t�5�	7|z�Ű�����$"O|���D͍B�b0�ւZ,<�M�q"O&ũ�؇m�|�$@�Ht��"O����cx#P!H��� t%{q"O�P�է�)V1�C"0����"O
�!�O:A5N�L��A ��d�<�ERZo��e��)@(<�`�b�<����2ѦA�gȁ;N/�d�E�F^�<����-Y0�����EH�öM`�<Iw�Yw� �
1��Z����d�[�<ّ�Z�j���&0�b7i~�<ID6
����DEɤ
��q㦝z�<yE;/�T�i�$��}Ԩ�I�E�]�<q%kL&Jcց�Y�L����[D�<�"
�4"X�Yb�Oӄ����c�u�<��=tļZe��>p�I�[X�<A̫Yx�5���/k�M��*V�<�O�0"��]�&��eHAi7!�T�<���� 4�ݠE̡N��5��F�<�ShE�n_�
%�6
|�{d�k�<qюD��D����\�F�:�'�d�<1 ����9�X4�bС���k�'Q?
�)I(=�`ЪL�
aPz���=D����Ȳ�|9�4
�6+�9�$�;D�PK��<�"|s¤ƴ$�x�@d�?D�@r�gP�qUr4$�`������;D�	�f��`�)�(J���15F;D�h h�W>p�+S+O���y4�:D���)��
m�&�ÀYU�|��h;D�̘�oC>��ӕ�^���h��&D��y�.L�w��S,-��1Ҭ&D�� @�CGΒ>���T�G-i��"O$͂���z5���H9�"O�9��U1GS<|��`�7i��q�"O� ���Ha��K֏��}	�4k%"O����:3�H����"����p"O��"R>C���x#�!Dʎ���"O� A4iɱ��=�u#�f���H�"OLt���M"dy�A��hP!�h%!�"Ob`�w�@&�$ �5��5Z8����"O��c�/�.�bH;�/�!S�`bP"O�q*��,q�`Ccn�LCPI�"OQ�U'�,#��(�!��G��v"OT��TdŲM���r0��B��[�"O$)�3���q��,y�@��pC��u"O��`�#|b��/��N�Xp"OT�j&/G)5��a$NT�$h�j�"OD�� nȥYT���r�Y�k!�t�"ONe�+�#)<�1� .<�8��"O֨���Jш�����T怢4"Ov���$މ?���[�$O�,m��"O���t�fj�4�a�J8�hd"�"O�K�^�o
�ͫ��HUu���"O:�b$�ƥXC	ԅ s|�+�"O�	���Ul�)��G�MpL0�"O���B�2�b%���Ū]T�ّ"O��Ê�h��zeʑ�qW�Ū'"O��+'�F�t?�p��k��I�Z�;f"O�`����f�(�k�'ОZ7����"O~$H�-ÒFN��fD2Y;t��"O�*bgZ�#eb�S���s�:��"O0equ	Ku��(��P�,�� �"O"�����(�Eт	[��"O� '/\���90tA[9$yʔ�V"O�3��%[�� C@�g`���"OE���C-h�183*;_�1��"O�Lj�n�:��x�5�e?�U�""O��Ȳ�K�yL�
I��5ȸy�"O�)x'Fɛ`R\�h���V5����"O�X�1�N�\���B��G>�	�B"O� �r!ؤ���nt�"O��Q��F��y��

VP�!�"O��YbO]�|,��;�G�]8��Zp"O��pB/rC*c@�j�||��"O�YeIY0C��lx����$<�c�"O��0��KU��U��)1�\+"OmY�^᠔��хh��1�"O�.-�>��ӯ�OP:u"����Py"�ց-�j����
E�b�Q��KZ�<I�-s}�}�D�]��p���V�<�6CQ�;l�У��+~6�0�jYi�<i�g]�K{F�X���[��-Z�<� L= �lQcs#��:���ѵlXQ�<�0(#b8�X��aX $ìzr�_T�<�A,�K���Ҡ]�) �Y6j�P�<��F��Px�y!M�Y`��N�M�<Y�͆M��$��U���+��1D���s�F��ˢ�Ӭj�ȘR�a5D��� ުw� 񂄍Тi���kw�6D�:�g�vhLŘe���fc� ��9D���Ɔ��~�C�'s�Uː���yr�%�:T�T �&S,B�@�W�yr���V]ա3�,_� )�Ŏ�y�U1�6��f�*{����G�7�y�*�dxi��9ykv���M �y
� �}�r�32L~)�+��+9֩s�"O�X�eaC�*S������-J.t�!W"O8iXt]�R�2�R�)�����ac"O�0��DP����"o_L���"O�Q�F�/J�f)S'�4Lvh�if"O�y���D��|���T#qj�أ"Oh� &��jU�:A�� Ag�x��"O���E��}�# �2G�*�B�"O�+V�$ ����3��d�`"O���I|"p�5M$1�*d(T"OV���� )��1��)�*��"O�I ����.�2 +S�V��Yx4"O.|S!�E+b���1ʋq�t�*5"O6�k�ُ,�F@�R/D�&����"O|ԙSlO�oB9aڅ8�ZP)�"O�JTIU�@�����`F�p-�y�3"O����ھ�\���aC�(/0��&"Olժ�ӾQ���2��],��H�"Opd��@�l�%)� ��!:��"O�j��@g�`�ѧ���QPz�#�"O�E7��Ba�	!�Ղ����hL!�ğ&?צ�w�Tz��	d�S�`�!�Ro�^���A�=d�p9SaO?.I!�$֑"���A�Y2)ZU���Q$?!�D@=l�d��R.. ���cD�!X�!�մ�H����W�f�r�ā=S�!�Da4YٵBW�C�2���d
<�!�Ĕ��0�-��0����}!�ߦ ��� gɑ!��XD��2!�!��+-�����=$o�D�t&�:�!�$�t�j���&K>cM�!���@��!�:pk���SK��H��#��<!X!��RA�$��S�PM�T����-y%!�D�C/
�@	�-!�H��/!�d��B�pZ"JՕ:�k��(j!�Ĉw �����\�|@��P?$!�;}Rp	��>8-��SEN�T�!�ď<^��1�ȟR*v�y�C��%[!�d� b;��B��8.1b��O�!��1H8)�b ��rWk�59!�ڴv/\]qE�F�!ZR�qEH[�I1!򤂟g�A��L> A�Hz2g��3<!��>�Z�����<=0�ك��}4!�$-2l��Fk�$,��	��'!�[$�\�p#״<�xB�Е)!��g���آhƞ7�4ٱ�D
!�$�4Xޠ�Z�M�j޸��"ə'�!��C�3�Tx���+���v`�	,u!�$VXQp ��ER�I~�R� �]!�'Dz�9�C͕ NK�.�>o�!��	X�y�T���$l�7-�6.�!�dK�V�^ࡢ�O t�~��W��1c���Q2%����G*� 	�y�ƍ�K�\h!��Q��`)��y2ɐ�a[4aR6J��F�vQ�����y�$]�vu��1Oq��j�5�y�E��9���c΀�Ha��⓭̲�y��~�4-�K;O��T��y�X�dfDyh��+�R�+$��y�)X�T���H� �+�
�yRaTv���n�a����oܱ�yRV4�2�Z7	�V��%*�yB.ѝC*�;��ǊK�hA D@I8�y�Ő�..��
)q������\��y
� ��3�ˁ',�|��T�6��3R"O:�20���)��H�#��/�
�"O�;��>.0,Д
�D`r�QP"O$	)��,0r��
l��(G"O��Rq�Yte�e��!Zv��Zs"Ov����F>Ґ� ��Y���1"OB�Y��M�?�2�;B(G;|�ȥˑ"Ot���n�Y�T[���L���5"O�١�� �*�U&"+�vh!#"O���fQ!�%Ҏ:��ܺ�"O �z���;X\^U
c�T�d����"O��zq�!��U���M!p�*y#�"O^�[�� vv ��l�b "O"��VKC�_�Dp�2�K�Y�}:�"O���G!CF*``&lN�&6�� "O<��mBi���딵 ���v"O44)C�w��9s�0���C"ON�AP-A0{^�8�S��xMA�"O(1a %��l�Y`-���D$b"O�p�%o:��Qe̝�n�%qd"O��� �6y&\Y�1��#��4"ORA+�!9�୍�Kj���"O��R�&O0מ`�u��!Q�F�@�"O�q�b��dx�PBʨ)��Ht"O��k�	E�8�<�B���9wԆY�"Ob\R��Pl� 5%��^)�"O����":,xH����5f���"Oz��f�Z�~���&��j�b2"O�P�"��t���@��U�I���"O�	�ĆWdI[Ч�	`1tX�"O:5���J64���E-|�
�"Oj`Ñ�ٛO�~m��E8���	�"O2��Ȕ)��i;�jJ�{��2�"O���"CB	"�U���_M�¸ s"O2 
���TM��p�_<)�H�&"O��A��wla����>�@dc�"O��¤,J9{�Ta /N�mn�e"O�E;V��R�,-ђ��eHL�ڣ"O��b���AK���N˨6.�a"O �z���i�t�W-�}��l�	�'0��j 
'"I�0��k�D�V1 	�'PR1O<I.�۷�������'��؋ÃC�y���C����$��'by[��� ��y"���8�2�'H~}�r�>z�����'V!x��'fl��}/����J�G��p�'�Z��dF�c����!K�;�L��'�ƹ���ڟ?}H�"�9Lp��Clli22E�#�Y�����*(�9�ȓ<@H���;#<����@=k~�U�ȓ<z`ј4@"���4�Q5Bb��ȓ4�������7~�&�ᆢM*?��هȓ	�Z)���$H�Ѫ�z�4��q:�-��aH�h"��b���-Ņ�K��1��N�F�{����p��qɦ��Ug�?`�]v.р��Ԇ�Lr��q%O��IZ��G&ZO�цȓO�F+�/E��¢%D� ���ȓ~Z
(%`�:ak(!��#[SX⑆�5�`qp�++ʹ��j�	�:��~v<�"���j�t��!C�X���ȓL�鲖-�-d� �va������'�.��6S�5
Mi�^�`����ȓ1b�EJ�'JX����P�|��S�? �I�q��0XX�QE5lL���"OX+��ւ0�Q�BʱpiL�""O��e�O�8�|��N�{��A�"O�	�p%�
�b@��o��`-.� �"O4aZ��A0L���mF-_ ={"O�H���5��"��%��uh�"O��Q![�b�ܰ�UJY)b|�9�W"O���&����p0�IY(5mX�"O�=��+��TX萦�Vtcj��"O:1�f�-��Y(�'a��z�"O�,�aN/r�H!��ՙb�B �"O�lpvjE� `��pq́�|<:l��"Op���ِ[7��i��4e��q"O8���L�7Ϙ���mJ(<�^�ҥ"Of�y� �4��,hcmW�<���"O�����U�^$b��ј /nt�1"O ����T@�PY�F֛m�<��"O4��)��>U3��C����iD"O�%{훏=J�����d�s"O��@��(OB!�G&ȚH�B�"O�Y۴�A���t'Q�~�Ȓ�"OB�i�nR5v�"da�*/��諒"OZD�%X���@��d�p���"O�ȸrm��9?� ����3"|l��G"O�ȉ�ňu��Ԭ�1�"Oj0�A��0oS�A��A|�4*�"O�����)�
#FL�.�.�S"O�d���?�jq��Ŋ�M��tK�"O��	#N�o��a&5yb�R�"O<��/�jlag>)x�Y�"O��gm�t�0&\�J�F��"O��J4��X�"4�$��t��!#�"O,̻Q	;TRL$G>`ؼ��D"O�m�U�ԓ��5
�Ě�?r.�!"O���6��lԮ�+�$?��"OB}���Q�mm.|q6F�C��9A"O|��d��{٘�C��R�R�Z%B�"O�d۴A^�K�q"G� �r|�"Om��6���"������8�"O�%�G�9"�^��W-��N���B�"O�р��O��0�T�T��"O~l#����$�j� �P gςD��"OT�0�(E�r%z�Ȱ,�/Q��{�"O>����PT�ʤ��"F|��"O8d"�bJ�h�*�V$R#�$
"O���0�. �4�#d%�38����r"O�<��A;���:"̙`��Y"OBȑ0`�7/����d���)�"OB�C#N�^���֧S�4Ő�"Oh���
�ۊ(0��w���"O~�Q"$4~TY�Q�]�� :�"O�l����?L�ģfM�f�~��"O�Y�L�=5'h|0�,ճ4VH�T"Oj,)��_�@�h!�U��7>���"O���@}:�P��R4��9�"O�}Q�\3-��}C���S�E�$"Ol�H�VFLp��Κ+
�#"OZ1j�%��qXX�0ЏN�l� �"O�x ��I�"ۆOL܈�5"O( ��	ӷ!���� �O*��Q��"O&�pW�H�w�C��k��RC"O�$�V	^��,�q'X7Β�9�"OT��`����Ԓ����x�6E"O�p��i�hÀl�$��$/@P$s"O� (K�äy	�%��W�`:l�I�"O2�SԮɉ*�X�X@`�.9�<�"O�T�B�B^���1勨[*�IpT"O,ȥ�@�JZYB�uh 1R"O�EiTH�3c4��aaB#M�%�`"O��;��/C��,��j�08J�`1U"O�tJ�흠|�j��Ɇ=�Qʰ"O�YCgȤl�|	P�MRB��@�"O<�@U�����O�T��U"ONTD(��f�`pB��P�I��*b"OA��*�O
1�+I	�D"�"Oz��p�Ӧx�R8���T*\���"O��O��1����Ôx:��"O����-Oz�`�fb�!9v4c�"OȄ;&/�h�F��"쁍{ �y�"O�+�ȉY�\`rT�3\X���"O��'��?	�!1aBP�0��<:&"O������a���BG�[��I�"O6)s׀/<@��b��|�~@��"O~�4o�<��"@�o����"O�L��W�q&�\..��%��"O
�+��ո/g$K,��V���"O�у��
�P�ؐ3���NuH%"O~��0#�0�(l@��Z@p�,��"OrL�N�Ao 0��g͊D��R"O`�	F�&(� t�D;��@b�"O|EIR�O!/�(Q�p�Ȩ�y�F"O�U�&%O� ՌE�'C!�=1�"OH�2U�]�u�2�	�Ş��D��"O����X�4�l���$�& �"O�	�2i@�Vqf����6�@ih�"O`L�v@�8����*\@�S�"O�!f�I�"tKߩ\�� 4"Onl�ˎ�^��j�'Bd1�"O�=��K]`ae�1(-��"O�D����+)����cĦi�P�rD"O.!	���`��Qb0 ن����"O@�1��&!XeB�� ��Aq�"OV49�;��Q� Ba�}�f"OP-)�L��N�F�E��AD����"Oޅ	��D�o�T̹�f�@����"O���A�4c��hj���?n�X�"O�)c��:A�x[��M�W$l�"O�e�X��L��#2*m`�"Oh�Bq��1iKʰ`R�#qU��"T"OX��L�j�ʔ�t�\�PT��S5"O����+U?�vd�T���c��J�"O�4��?W��2�mݮy7��j "O�)A$�&),.hra�G&�(M��"OFTZ��(NSx�a�����JQ"Oڥ��j
z�|���E�U����Q"O�P�(~�[�V�m�:I�"O��%���
` �A�kd�1��"OfajĤB�~��Q������[g"O�p�b��b��X'h�c�.��f"O�16�W(3q���a�n%\9b�"O:\A�.ɹkPޑ��A &,r"}bd"O�Th0&�V�h� �'1`z��"O�� �� ��pBs��W��U�6"O�-����=F��n��fʸ�$"O�$�歋/R��ؓC�~��B"O�`g�&��y!��/8n���"O>��R��+���X#�VY|��"O2���"�7��)�6��65l%1�"O� ��"���1��a`#�5Mvd��"O��и����p�A.%����"Ob�a�d�R�պeL�*�5�0"O�`�Qlˠ&��ps�X�����"OrTk$���=����f��[�D2��۟��&Ҭ_s����r,�Űw�W�nQ��S�!��?�]�P2H>����I�6@��iS�U$#���XE�=���Q��(h.d �!잙V�8�QFS��II�7@�{S/Q��*\c���e�'M*iI���?I�����i�����紴{��	R\�����O��Op�d9������m�yI�!SgFiu�d�C;�O��m�ԟ�n� Z�hd$D=�y�jM6xۼ �V�i��tbc��ĸ<y,����Ob7-
"s�h�OO="���&�(\�丰a:E�ph��OD�'��<�aDׂ3�`D�"K {�"(H��Ϧ�������IT7Llq���3�H�kl��x���:�\`�E/ :ݛ6/��?a�����'�?7�@8{�H�E 1V�Tٱ�â@����O���(�S��(T�J��~B�\Y�$X)Z�<Y�id�6m)�SϺ+��:oM
1j ��84����L��I�s2��ڴ�?����?IO>��o���`�)��k�,����Qc�����۠�5#�O�1PUke=p+MD=x<�@v}��O�o����2��xb�7'Q����"�ype�`�Ԁg6��>/D���OXx���	���'�����ڗ�~!'щ]��y�5n*$� 0ףԠ|8�`�Y/#��� oӄ7-�Ǧ]�<��?ݕ'�,-sr�F),k�iæ�u⎍c��U�����'m"�'ɧ�4�'zE�.O@��)��n׌�*��dc� ���'�� �ir\��;��C�~���I����t�ju���p�����.\��i��(0��P�z��E�S�>�⑁�N��@��h�S���գ,�>�����%bۄB^��~�A%�S�O|�An�W��y���N35���(�'�x6_צ�'�J�K�f����.�)� w�h�3z���We�33���?��o5ԙ���ʊ6Z�I��x�O����D��w^�Ԛ� ͟�JT����H�N�d`Z�.Գ*yj��U��ŀ �J���Ϋhj@���HO�����'A��u�B�$�~�AA&<�����/	4�Dए5n"�4�|"=��MI�(���/p�<,���s8��Xش.���i;��A�[�����敺z���'���ĩ>q(O���<����e� `�4+������T��z�iT�Q�"�x��'��	>Tv9�!&Xk�61�@$P=�7�F�PW0��Q�U>?x�)��̄�H-.��%��r���¤�}Ӏ�P!�'�op�2�$=���2WWM�tE��'�
j�V��T������Oy�'��	�M��4�f)�7�X�Wh�����{Ӝ�,���6M��"��+���7���׊�N��&�ȅ퉂w�� p   �   �  �  �    B$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�U曞@�VM�P������@��P_`���'4r�'d�|J?��f�s^hy�&A�x������ b�8�`XTv�|2���,�
�*��ڹz7"a��iRȖ:[�Fi��	�[ڀ3�F�\l����S�
��0ɂ��O��d�O:�d�<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&��|�����$��::�i�V�%C���e�Ԋ!�lK��O4�$�O��d9��~r"&F�L����� �45`� ��A%h�d��o�&=���1���Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�Y�P�{ � T�>�@� D�(1! " ��Eɵk��<�s�j �M{��$�~��A�(���4 ��7�*��2��y>���=���O>˓ I��"��ߣo��u�)9?Ԡ��F��r����y � ыU6��ȓ~�p�k%��^��1� �
$F��ȓN�� ��啦 jN=H�Aއl�І������(����� #zy�q��K!�2�"MF�����X���KV�w<�%2�M_�I��$�OD���B<�����J��`9���)�!���r�¹�P�D*/���2!�ah!���#S_l$�f��dQ�ݒ��߂*L!��F
�L w	�zE���'�@�H�x��#���P�P��Sap��M:L-���J`eEx�O`��'=�)� (仃'یBx��"���6�˰"O�q@�	��@�aKb�1h�Lm�"OaP����`��\���3��"O���lr��-�3|�z)�u"O��vJS�-��H+A��usp	A��>i��)��1j�L�B��ΥjՈ��1��+���'*T��d�'7B�|J~�A��99�p��G�fp�3�C
Q�<Y@��d�f�B;R�&D�S"ML�<�#ۼ|����#��(���H�<)�MםB���5
�=bxD����G�<1�Ç�;i��aڡb`�Ց��^ܓO���u(�O�=�S¤�BHC�e �s�۟�&��)�gy"lG",*Ȼfc�7hs����)���y�Q^�H��0��#�$��y��O��z�1�
��} ���qAϬ�y(RC��U�?A���I2F��Pxb�)�Ql��\�pH�Ĩґ+��F}Ҁ�:�h��=a0�A>�R��g�*� �ȝӟp�	lX����O�N����ql �Y�b@��;D��SvA�zb2��Kߺ�
T��=D� 9`�_�#X=R�H�8����'j8D�8���_���K��X�Y�(�RT�5O�DyR�G:nJ9XC�+����W�L��~2'��O�)�Oj���>i#�\��:�b��Ǒ8���k6`�V�<�fM�iH��&k�T5P�Gi�<y��
i���uA�&/<�� �Qy�<)��8
;�9$N�Y½�eQZ�<�O�3��2&
�ڵ��QP���k���O$�9j`&15ʱp%a�m����I�h��������v�)�i	0�
�ː���3^�M��LGk+!��;m&yBQ͓�`���k��H!�d�,PD
���/�|��Aɂv%!�$
ZO�9eD�J�΍�s
B�!�$PGS.]*��;��xH�jqO��D~2o�:�?)�O	�s�  ��ڙpmr���[��R�|�����I8)a�<�7.G3@O�t[�/�Y�C�P�2��¨-��X�΅=g�B�I�x��u��
�&%^��#�
�T�vB��*H��!(9�`"E�^�hB�ɛ0��!�@��� h�BD�H2�Q�'7�-A���L"<�X�a!���C���&3���I֟P����#��� ���9�h��(�+T�B�I�-m^��qJ\�{戔s�/	�ZB�ɸT]&� �Q��\�Ї��LUXB䉌v�>���Ã6Lh8��l�p�J��D�q�'���c��ƙ��%P!�ۢ��(q�'�0�K��4�����O��[�$%h����$u��	��[�$`���&�A� � Gt�$5.]�t?F�ȓ|�@9�e�-Dy���L$A�bф�b+����`�����lr�ȓp��$0�&��i�w�>�ܴ�O� Dz��4&ɖyy�p����>'˸@
�����	��š�O��$+����m�����.��"��b�L�yRD-k:i�4O�.0E(%l��y��X���놆�
}\yQD'˒�y�g�m}�p䃏�z.*)�����y���==u��AK&q��ih GȊ��'*�#?�E����ܓ�L�hFa��]8��!�=�?AL>)�S���'(���Z#��hi,���f��MG!�	:��ѡp�Ĵ3&|���R*!�$D(7�习���@Jm:�A�Vv!�d��>�p�$ =J��9���+#�𤜠
�\+%�3y��D�G���m?\����
=��>q���^ j�`�v�Z{ج)!���?q��>� �8�G�?��L[�"�)b��""O,����s�����E�<��"O���QfFI�Ѝ��:{*�Z"O|��ä:/pCs��~����'B�<�ޯW5� S���2.�H3L�{?Q��Fe�����'N2]��`d\M�֨H�@�!qg����:D�(�GزV����j�+��E� �#D������;%���s�f�$.A�\I®!D�TK�b�+0���딡!v(I"�>D���hB��(��EƬ8�<�!u� }"�4�S��L�����J�/vJY[3D͜<�q�OiIAI�O���3������8���Y��Y� ��������y��E���[�G��jP��!Ð��y"/��x�P)X�e�H�R!�Q�yJ^��qႨ��a �1бnD,�yBeܜyd�� ��*� ��@�C��'�*#?� �Ꟑ�g�J
�pt�2��4�>l�V��?!H>��S���DX�^�XCB�Q,�$2S�]�,�!��.�B��#$Z:a�*�w���W!�d��~�U
Cd�=H��e���v�!�DM�(������E,<�Vy�Cm�F��ā+M����G^
xL"6%".��$�>����X�s�, �W�W�}��5[����?9���>I��� ��p�j�.c~��R�cGS�<��C<o�y ��w`R�+�J�<.�Qھ�Jć!�b!�*E�<�2 �gm~�`Fĝ`��;#d�\8�H����-�L�ە��> �ݡ�m�F���I����\��Y}��Y�5�آ����9��9{����yH��E(
%Q����4-�Ա��yB���J�`��)�$4RJI	����yB�[�g�X2'm&t�H8�hO;�y2�6Rzp��Ag�@بCoA:��I��HO�$�zwΚ�����$}}�=��>��֑�?y���S��q��yC��1S��Vi��C�	�N�NhT�X9T30��Q�ˣ8�bC�ɆP�ɩ�X�"`n�(�+�%tB�I���B�aҀ`
t��E�I�"B�et@�@#� ����G�U��X���<I�� cNxԙ�	J���:U�C�4���%���O>���M1��%?|8�a4�������E����s�Iy�G5�&m��[�>1�5C�D�Xu�QF�"��ȓJ8���J}R8�3D˺%����~��m�5L[�\��`6���҂�#�#<J8G���
,�(���:F�x��Rɨ�$�O0��:r=��@�շ9��Q{�M�@�!��]1 ���q�+�9`E>컕k�NK!�Ev�iP&�%Բu�a@Gb,!�_�vpi�CV=��1�i�-%��xR1� ��M�pk��<M24⃋��\�X��$�"Fx�OL��'���9L�r�&��v84��H��$�C��$q��
Ѩ�9#fԨ�j@>1C��"h��E��/לA�����%J+�B�	Lb9�ÆȀ	#8t�V"�x��C�	�q�z0�e��#�|5oZ!P��'�"=�z����2cj�Ј7�ʕ�F$�R������OH��-��	V,MQb�ɍ�3�24A��5�y��٤#�4��#w�H�jA�Ҕ�yB%A`�V%�q�Зo*���
��yb*K$���΋�R����m���yr�B���\C��#K��$C5����'�l"?�rʟ�˳��8D~�� E�MF8��O��?	K>��S��򤗗g��AB�˾`{"(��Iս3�!��  1��e@u��8���H���@"OԌ�e�^�2��KE���+����"O�Q2+_�F	f� �H�#�ܤJ�
OV�k�3+��2@@��8��e�����O��H��S+�~ ���ͼHqh��v��!+Fȵ����?	�	<t!�̇�: �A ���E�4��ȓF��dՋİt���Õ���q�����$���7(ܣ�����'�
@����+O�UQ�*�Qo���r܎- � ��I�(OD)Q�*�)>��y�5�Y>}~����O�rb�i>}�I���'\���צ�1�P��-P}R���''�e�T�;n�z��Oչcb���'c����f>w�j	����X3�1�'x�`�􇎋@.��%�8f�t	�''4� �=/z�B�.�3W�>�N�h����)&U
n(z��N<3A��IK����|�����?AL>%?��S�T��bP��N��@���?D�$�f���T�b9ص́�?U4Aa��>D�hơ��b���'#˷Q��v>D�V٘ ��) E�s���	�Z��y��Y��r㨚(g/ tȱH���'��#?�0G�ן��$DٚR+��3�Y�&��D��?�M>��S���=4.� �偙�s�0%�r�X�E�!��<A��#wA�9��h3��be!�S�c�%�%Y�v� ԩؓG-!�d.]T��4�hr�`M$���Ȼ.������-7VP�1�D�_���䑞u��>	sg-��"�u�2��!���7똰�?)����>qV��
&�(l'��#iv�r�jc�<��aA S5Z�颥�\�>��q�_�<�aP� �n@�6��$����K[�<�C�x=\H�&�P��0jN{8����dF�q��)�7G�b*����L�/����n���ϟ(�IC}-'hpZ�
(!�[*C����yBg�0�,A��R8&�H����$�y2�Еf��͛���+"P>%�!�\��y2��:�ɥ��lr�@p�ۥ�y��Y�"�����m�+Ro�� ��3��	?�HO�2��4�S:\�ҁ�&$s�4:1�>�0�ϵ�?i����S��/�ё��~\ޠp��Rw��B䉝2�8d[0΄ifzR��bM�B�	�p��a���)C�j���k�Am�C�2i��5mޡoX�Q�gŏfKdB�	4%�]H&/��IDT( !D�hJ���r���E-/��8{���#vî*T�ç!ͤj1��d>��O>�|��������pL�Vc�=�y�ȓbTȁ��N����q���T�O��#*`88soK�F-|��g�1m�,�ȓ��e.؍\�nMb!B+=L�a�rt�G���;jd�!�V��e:�=��r�D�Td�]�8<	VX+8�*\��j�/XE4���O������t}�DÐ�:z��!���M�!�$D�g�����?q�8;�-g�!�d�U��i[ �F&�ƌ"�m߬b�!��ں�Kg\;� �6Ώz��x��"ʓ{j�P�S��)��a�D�5W���E��Fx�O�B�'��Ɉ8�
B0���!�dJ��g�JC�ɪ�AH��ep���GKǋG�.C�<7<D���>�Ȱ�7!B.Y��B�	�i*���M�Rf����şz��B�	RYРs��P�P�wiɸ ���'�^#=��얶g��m9T�X�	�.��@cQ�D�7� ���O��O�OW�s$��)b�����?&��'G�P�&�"���a��,A���3��� �]ytG[�7���V��To�i�v"O4P�P!M{�h`���h_���F"O6I��*�<6���냁�E^z�`��d]�'�fX"��V���R��T�l�%���Jb�vje�'��'���Y����,J�,�@���ܖ.X����*D�� �mδ��S�Z�65�'D�@c�b�*դ�%��Mʬ*p�#D�|���A�,s�$Zu��k�֙�'�+������v���IcN:9�T��m�3XQ�$�@F0ڧH��Y�)Z�Xl���J�J���'���'�~���$j��`9�c��z�0	�'aRX��e��$��Hi��F-Y��1R�'y�Y���%}�DI U�?_h|P	�'�f�
&��F.�]9T�P�Z6�9�
�Q�Q�{��s�u���"i2re&�i�'m�Y��h���O��V\�ؐ���%R�t�>o^c4c�-~(�k��OpTR��j�g≽[т�H��F�w�� ��@��Y�v+�6.�`j�'R&�A��4�3�$�_ Y�%F8�$)Zi\�|��	y~�jҸ�?ͧ�HOL0D*�a���8bH��Ft�4"O��vH��29�g&�\2����>���i>���_}b��h`�hrV@O �zH�m^�I���
������䟀'��O�\�("mV�{�DՒ��ז2��r�N����4OP�{[��X��'�d-P��ҽWh�a��s�h��Eʟa��]��8�J$�'��	��i��?ҙz&��
L�2�m���?	��hO�c��(6�l<�|��a[9��Bi9D��4 X;��sE\���Q��`9�	��M����'k�����-`d��BW��Dӧ�V4=���'1�'��Y��!�{Q@�Y�'�<l{BJ:D�h����355�����	WB([% ,D�(B���i*lAT����iiG�/D�������L�Y��T�&3ȕ���.�� rFD=�<���`��C��1���LdQ�(��#<ڧ%�M ���]�Dmz� ���1)A�'o��'�ڕ�P�H
�x4�n�@Й
�'P���j.X�F�B
�{�@���'�b�Z�m�O��m;�I��/����'�����t���� 8�(�Ǔ_Q�D ��!\<��d�m`���Sͮ���)��|����?y�O ���h�-eڴ����L�1&"O0��Ӥ� {v�q��øq)e(�"O� �2͛1���րQ�(�4x�"O@����$GM�[��[/u�|��"Ox��e߭lh�QP.G��p("U�>QT�)�S ��M�*�h�´���=����wb/}r���z��'ɧ�'>/�J� �7=~th�O*�,��zLi��L�j�x`�u�P3�D�ȓ�0��1eӘiA���g�?�\��_��*���K�����+r>1��M�BuҦ�"R<f��clм"6܍�=���I����$�<C�!�JE}��J��"VzBL�Id�I�"|�'���vDL@�pPq���Z���K�'|X�顬�.JM�)���E�R-����'��H�B�	 P*�B�K	�BY4��	�'FŃp��3L��m�$�B�:��
�'\@@��ӻ+6�Q	A�ۡI�0�q�{�'W��9�'_�2�����7$zj�)�K>pQ ��5�'��'ߠ��2*(���lY!zc�0
�'�\k�ǖ�pL:L����wt2MB	�'R�7�Ļ5iʠ �l��}8@��'��X�_9�T�ʡ�F�!���ǓQ� ���V�����(D'�p|Ȣ�3D�����  �    �  �  *  y  �"  �(  P*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms��a?Aab��jD�O�,P���$�0y�x�����A��j�w��}�n�W�R��&R~��YBd�*���$� y�~`#_|X, ��o��L�#hZ�i$��`N:�`�O��t��XF{b� �v5��-��.s��c"ճ�~�Ƹ�R��!dH���J���7�ybf�9b��a��Ƿ��P�F&�?!D�V��|�¬�,�`sgb�i?�"�%̓@_����duP2��%�y��K%i�i�J�PLQ�ALR�>T�D��f?i�f��."�O=b@�V�DS ?G������_�h�n��0?I��Iڂ�8�L=*���ؑ�]�s�z�*5�X�L!LԢ@K��=)\9��_��0=�F�]�"�vT�YI��I!G�&\5ўԡD�U���T��*]�QHh������]�p�hQYB�G"{UlՊ7�#D��ٴ
L�K䱱"�D �2-94J�O@��@Bδ �)ۂc�T�ض�O���`ӣƠP��/0�jD��L-D�ȹĬ��s��+�G�����-��k�ڈ;��O���b�/O���'^�~(�<A'IL<{.�Y$�j��ط@Hvx��ٵD@&T�D�2��A�!,V9H��Fe�r�G���D�f��$� �`V"�q���S�˓I4�yb����l�V�Ha� �"�TA��`M���#c)��5{��!�L�����ȁ�g���ȓ�rP�5�ڛEC��!dO�	&���	%}(�X6 @b��a��Y�;���)��40V�e
�Rw|��&�C������4�|���62�V�h�����8@q�'`���I.�5��é|�D�ۺ��'�J�(���j���ɕ	��s:}@�S^�}Aw�ܟ2ܠ���� 9�
7n4N?���		P�8	����P�v@��l��VCY�-��Q��[n E{ @@6�QTbóX�4� �Ɇ�~2�J,")��"@a�"� IZ!L�-�y�	]5'�ҝ@��(�Ҽ��"���?q�(�$^����*Ż(l(��Ue?�r�K�}`k1��Pd(��f#��y��{�ir4�
hjR\���=���5
�v?Q���f��O��@Q�$��@��r&�d�f�#���1�}"���$q�Ț� �����G)~��%*������H�_HΌq���(z�bi�C�'��4" ��k��)�(����EI��$��͈Ȳ�Œ8'%
%K2#4U���0k2�� ���������O�]f!� �a|���W�;M،i[��IW�#�^% �҆ɐ��J��v���~���IXFr�8�Q�)?
@��l�E\!�dٛ'i�*�KCRi:���ͶZa�x��S��~��f(6�)��ii@.%�I�{8�ԏL�$�����2)B��"!i�d�����Ed��°��Y��1�0�+T
�YFB�=,�~����)�n����3�Б���I3j��rd�6ў,��*T$n�hЈ�!]� �6����ȓ$�Z��� bBE�&��d���$D��7=:N�X��M3��J�i�	��̞^4�2P��6�´���S�'QƀRp��;R���P'F)H�.!��'��4���R01�g� xt|�8�*G��x�#����o�Y��gQ1O�٪D��:R\��f�/V��4�""O�b�@�TY6�G/\�]� ��"O:P��F��'j1���20���"OR��!�CY:��-ƆO}�<`V"O�����+]�Yr�͝�]�5;`"O��C��,���R!�*v4�@"O���e����4���|V�\ۤ"O�P�#/I.��zU�y@�M�G"O��iҎef`�b��z�41ia"OL�P��
eڰ�B��>h�Hȡ"O<����&�&,�Co��`�����"O�aQ�ٮAf���ݞA�a��"Opy����L#��1BM�4%�U#"O�,�l�>p���$/^IwbA�c"O��؅��&Q�H�aM�>?�dr"O,aYgi'A-��BR�:=���Qg"O�����gH���S"ۼ#�H�5"O��@�#S��I�D�23��_�<�MG�:�m ��/x`�hq��W�<��hڜ&�|�3����"@p�"V�<!�o�?l��aV`��a�j�ծ�Q�<�uG�\W ��𩛔mY�iNTQ�<��l k�8u���֐<��%y�e�c�<A��DIU���'�s
ԡ#$JX�<���<�
�H�I�X��a��o�<��\�-7�!���>Uɀy��C�<�ŊҞ10h��> ��Z�j]�<'�H��z}�Ì%�� t�M�<Qe�9��@`r��5<xt؆"CH�<�QW9<ī�-�n)�Īs��\�<)r�Q��,K�� +���
3E�V�<1s�=f\�zu�7�Ig��m�<�uF/��|�4k�+22n�t�b�<�pbV�D���I�Dg��|;A�a�<�W��3��s�	�t��}ZG��h�<q��ƌ65.x���k��5r��K�<)s�
	�j���zP`C�<��h !�4Kfj,i5��ˡ�@_�<��;yFy�dϩ�l����S�<YÈPV%Y�@ͼg~9��OS�<�5BZ/Bf��{��Գq#�!���CQ�<I�i��9�X= �)B�z@0��Y�<p/D�'"ȍ'�%��cU�<�4��#m8d���K�jn:<{�I�<ɧ�
T	|}Х(īL��0�A�D�<Y�j9�p��q!��ܹ8R��h�<�q�W
��:��$^�ʙ�EF�a�<��e�,gV�l�����\XȔ��B�<1��ڦ"�䛱�ײ��=�Z��ȓ<��(�Ǧ��*<��.)a��E�ȓ-
�CF ѳ5a�c�Ο?q�����S�? ��@BC��B�a��c��h�"X�"O�a����4�@K�B���}��"O8�ā^!Of>p�3�C t 9Hp"O��G*B�zD�4!��$BY��"Op��A #+:�� ���$._�D�"O�9����8�Q�M�DE��j�'��*H�9�4�fEE�_�6P��'U��8D!WQ�\HQ�^nU+�'���1`��	h,㰭�Y��Ls	�'����͂�mϲd@@$C�V��r�'8��ʃ�ޒ;e���$�EO�>��'Q�H&d��b{�0�T�p˄�	�'s�PC�-!Nv�h���}�Y	�'��};'�@؅ic慭t�� ��'���s#�G���k�c,i��0��'�Nx�" O69J|��iׯn�^�K�'�l�z4�R�2L��` BH�pN0�'!:̩s ߷r
��3@�"|ծ|p�'Gmh��6�^�B#�x*�x�'�+o�61h (%�.!�U�V�/D�` f��L��0��8T�Y  N:D���� ԛH9��{� ݔ�����&D���M�mJP8�癢k���R��%D�t�%!Y�,@�i�v�X�9ž�Zc#D��V��Q0����o��P2�<k�d D�� S�@G�����Ֆ.^yȆM.D��A+�9Æ8��F$�>��`�&D���5̏�u[̑�Fj&2[4A$D�D'���+J��p��#g�2�1!-8D��+A�יఽ�T��_�m`�1D�|�t�;;8.<KAM��ۅ1D��p�B��JΊ���",)�<�e4D�|�*V�Ghn	�R� V�t|��(D�h�T�\��8R$����K�f5D�x*HѰp�u�@�b���W` D�j#���>p�C�D�|8���"D��� �I�q�M��Gn"<q��!D�4b�)ރ�f!���P2���j@m/D�4�P�Y�Q"P�2�O�!?,,��7D�t�J�!>T^+V��5T`�i�6D�<É�/�nhhuD�#B"��F�2D���I>���S3IC�	��4J��5D�<+��1i&�ɡ&l �L���E3D�tᦨ	{�``2
ϯ`?|�!"�1D��xR�^�����O���"s�?D���!!��m$�I�ɉn��B6�!D�`('�M�N��p#d����M�W�,T�pr�*�@����2hֺuؕ"OVaʰ��t�`��p
��=`"O(��LP$aVV�q��<]��"O�aJU�[�?�=��L֋xYv�bR"O����*,�,@��V�
_J��"O�x��k�X���"�l�n�Hq"O����+��"��vȶ�Pq"O���O�%��ՑD74�|9�"O0���x/)��O�2���J"O��c�m�ϢAc �H7'�2� "Or�y�̘�{NѨe&םUBB�k�"O|�
��%0�2� %	&@ȑ�"O���𩇡 G.<�&���t�"Oq@�I�l�\ �B��r���#"O�<�7�ɞm/ؘ�oƱP�%x"OH)H���@�Ne9.��sz����"OĔ� �ק�r�{�NS�Fx��&"O� �X��N�C�j��5��vq>��P"O��a]�- ��kN
*prmi5"O��f�/�X�	���2F�u:�"O�Ih��B<&�
��6`<ƒ�k�"O �r�Ā(�5��-T�G&��W"Oz0���ә/"l�L 3�Ģ"O�8v�s�NԺ��:����"O�A�&^�81h��t�ڏ��$�A"O�A��dY������GͰTy.�֎{���/B_X��J��!h�؀i�̋ ;���@�=D���I��xz$��:p����<D�HL��X����ؘ��=D�4�hC/VD�(��׾�\����1D���c�*����
	�N�[�,1D�p�T�N���l�e���Z�,,�e`2D��@�J�q��(`!+�z�<�&�1D��P��w��XD�.��0��*D�H�
��q -H%��I��;��)D���g� �?ab�i@E�S��}I�,(D�L��	�_��9�6#
��:D��)��˱H�Hd���D�RJ�S�'7D�S��=6Y���E>aT��'F!D�x"��ѐ�j�zjN�M�X��� D�3��A�z�$��%@�8���+0�1D����ջ:ڢ�B��wv�]�� 2D���	g	Ƒ�wj�1�#%%D���b`F�gyn$�fǋ�q�~	��I8D���T?���4(=�����8D�1�%U�{o���*�C�f�X"D�<�%2BW��"M ���K"D���eN�']*mBC�ðSx&��!�"D�<��X=Lu�d�򩀼-�"x �@!D�T��Hߺ�HT蜔W{4dB3+$D�����={�Y�"�P����!D� �r�¤��K&g�q4�a;SO#D�0�2�^����ĭX����ej%D�t�c�F�<*4�&�@��׉!�$��(>l�2�T�<[bI�.�!�ć(hЄj�-�t �S�!���[��y U���`��M�@!!��!#Lv�P�ǒ���D�c!�Č�J|8��_7����:{�!�䈸�h��򎊴 ?8\�[>�!�]+�:1"Q�I|%��*�+\1!��M�U��JE}	h;Eܭn!�Đ��x���~�B��E�Q!�$�_u>9��A'�H �&��!�DL�,Hi��f
�~ɨ��U��!�d]�����N	~ D ��%v!���������3^�L�Bp�	d!��-�}�ģƪR	��Y�J*D!��ҺsY�H:�'�
S�@��e�,V�!򤎿b��� B)C-�QY�D^%N�!�d��GG�p6�ͷ>�!�5^6wy!�M�-P�G�0k���4D�c!�D:/t�Ȱ�)�]�@U�c��S�!�	'�T���Ȱf��DI����#�!���}�$�2�"�t�`̹��1	l!�Ǜ.������ծC*�j$�\j!�#�$���n�q�*�qFe!�!�ēq�"���'��v�L,_�!�ǣy�$A��DK�X���fd�6�!�D��5h�q9�LY9i�m���Z�mN!򤐖q(�����c��	
"S2!�� ��YC%N�o�Ha$�_��-Z�"O
m�ǩr����cA,lF$�V"Ou� ��T�
��ͼB+�Q��"O8S�a�HoFMA'FF�$�<��"Ol<!��[4H� �g�'|g�|�G"O��qA�hS8g r@E��"O�`��F`��81����:;�M�e"O�y2kӜ%y�,�����u�S�y�L��0!v��-�,�xt�K(�y2�F$E��qeO%#�m��,S�yr'�)dH1���I�$�h�� �y�ĝ�*9�y���mn�Kw�Z �y�n�
s~Cbd�"j|X:N��y~"����
^t�=j���"�y�"\�������[�h��˻�yb�L�k<ܤ)��N!U�H�f��0�y"DՍ>�D���Z�i��4��N��y��*ֲ�r�j�b���� ���yR��0�p���m\7G�t��)	��y����44����ד��X��mP5�y"�R�
�ڡhӄ	z�24s���y�oY8NJ�aǠQ�_N��j�7�yB�˭7~)�Ώ
w(�����y�K�ml�@��L�Jxu���y2DT�%v�!����i+.�y2��>��Â��z�����H��ye	/l�t�D(F%$)��ē��y�,�aH5(4eJ"xp!Cgπ/�y�)�Vvx�n���8�q�[e�<YaD]!5�СG��eQ[��z�<)ƍ_$1x�]%�PL����Hs�<��`�*��Bg@?Y�S��g�<A���cĸa���)z�J�de�<Y�*��26D��N-5�P1F�Yf�<I����Vd�Q,C7����&l�<��͊X�@�q�P�;�,sÉFk�<����C�t�2䞅~�)K⢛�<��/@�R��|����LdB�*�*�f�<�!嗍i�L�Q����Y Ѣ�dZz�<Iqi%v�*T �K�8�r��Nt�<�s�QY�����/"2Mra��w�<��%�0S4�jf�0Ht�Bc��]�<�TŃ�[;TTA�Z�7_�i��i�r�<AB��5q��i��g\-K.n ���j�<�U����y���ڏ\��2#�M�<� m4���cM�Y/TAb��J�<)���/	z���F�'t�>����G�<9$�Ƃ�ph�#Q=��Έh�<oR�}1��镎�D/�I�Bmo�<���b�b�B[ .t샧f�k�<�&Nƴh`���"p�$��m�N�<A$�	�:��R�	C�]��� ��S�<9���2&ּ��k�>f ����a�t�<�@JVj-���!��j��(�U,LU�<���?���!�Ο3u ��w�CQ�<QF�Y0��`�O�tl�"��M�<����?Ճ��N���s���J�<�c��$�j�Y��;)�� 3�@�<B���q�y�VMA�6���"W�x�<��ME�'�j�뀮�0h.Hԛ��v�<Yr��r�D!�#�,J����g�<Q���)��4��l��Q��{���w�<u4
��ib�ʇ�72Z Qb��r�<Q�'P Y~`�&H>'r ���,v�<� 
(	�GɈe����M/T�ӥ"O<���CF7,��
�6\��A�"O��a�NS8V�j�s�H��/� �"O|j��"�%�?D'x�yc�A��y"m�L�X��4Rv2�dY5�y����� �`�)Lš�-��y�䍘��艕E��Q�tY$+��y��է=זѲR�L8:�p`�ā��y"'�.)&����9�`A��`X��yr	�<0�J�QC74�Hg���yb��ZLɸ�8)j�#�M��yr��C�8��c����9&#�$�y�@� ���m&�6��I]&�y�B
CE�I���M����k��ɟ�yr�X��	��*P���V��yB�I<B#�)��D�>U�n8V� ��yJ0� �86&ݶ~1��h����y���=äI(���oJą!Վ���y�#N�#��/Ċ`:���f@
�y�)�9U9�s�T�QHErD��y�o�>�4Ht����P��D�y���8M�5cnB et �H��y����
x(cAK����F��<�y�JK�,�B�˵�+���S+�y�IC�:m�[��ҫ �j�9�,� �y�D f�%�C��x��$�3(�
�yR+��	�	���O�h1�廇�T�y2B�T�\-��	ozT1�J�9�yB���Sj҄
eH�{�l=������y���5y.�A�u�΅c��%X���y���"
���1��Tm�FEc�$�'�y�	�>�x(P�OY�c�f��@"���y�߶[plْ� ��u9����yR)&?8�䙑��X��1�r ��y ��`��iK��M���1	��yb?�P�8p@�v6 	��)���y�`C$P�)Т/4�ZH���y"���'�<�襎Pc������y�ݙ��Q,U��A�#���\��F>l�Q�]�o�� �n׻�FĆ�#ڞ�˴%�Uk*�k��l�(��R�=���׆>p����H�%���ȓ$���+7�}�A+p ɐ�����%���>k�T(���^.�*q���jM	��ٚ 5��A�+-{����+����@�fYD��	�%'n渆ȓ1��ņ�(��h�I������)z����P@�#fD�<���ȓ7$���>z���0�Ɲ A� �ȓN@����M�'�6�C����$�te�ȓ�D+�L˓��\�D�V�4��ȓ0�hx#0��,QN\�'J��&�N���ҺRF�
^F��9mH<��5�H=(qcA�,���&Y��l��|����#�W��т��O/U��ل�E*Չ��N "��XB��èC@ P��o�6�aP肍Z���1�	I" ��-��}`���QiA�d^R ����t��i=0�
GaI>yLl��E�ʘ	(d��R�Iۧ#�.�U������ȓ�~�۷�^0z�m�Q�F±�ȓ^z���"I�q���c0d��Y��ȓ��@A��Ch;aJ�5�؇�l�|�@�(���W�G���m��S�? �T�W�G�2m�p�K\�vp�R"O��Ô��*?4�<r%��
�x8�"O��SRk��
.A�Af
�M��i"O�,��_M�vL[d�M�PQZX[#"O~�򢏂	X�(8��ċ=o4Yj�"O��P����B����3Ȍh�"O�<�Ǥ�	�F �գ=�N��"OTM�ğ�>\�1y��Z	�,�"Ob,�ҁKZd� ��@�2>}h ��"O���f���<��
۝OxUp�"OD�fm�v�F�����e�� �"O�}� %�6,a��3[RV-9e"O�(�F���{��(� �J�ɲ�"O ��`�  ��   �	  B  K  U  1'  ?0  ;  "F  0Q  +\  h  Gs    H�  �  ��  &�  ��  /�  ��  .�  r�  ��  ��  ?�  ��  ��  2�  v�  ��   a � * � ! �' �- 4 U: �@ "G xM 1T �Z :a �j js �y � �� � M� �� ͥ �  x�y�C˸��%�RO5d��p��'l��ɂBy��@0�'�F��A��|�^{���OM4ب�h�e���N*E�M��_/U�LD ���Uq������}�:�ݠtX��ӤA:����xr	2a� K��E�#rޒ�@�,���:�h�?X�r��qJ�|a�$�\w����O�d6�ͯx�.�y����]����
&r�mà�C�v�bP�	;� �����s��Yc�45�������?����?���k�<�q'�An�XU���Hd�ar���?��?q-O�˓���O�EQ��"$F�h�f��9=�X��1G�O\�D-�$�Oh��R)����<)0�ǧ0T�	�3*»zGBI����S�<�DF�43�H��6E<J�R�o�П��Č>����3LK�
 x�O� C�ո(��=���O������d��};�79��(
Q�'���'���'P��'����TK_��%�`�͂���Q�h�8F�2!s�L�m��Ms"]�D�ܴv�ľi��� TȚ/�]���0�+�	����dP��ȟ ɲD�L(V�ي�k�$%
y���'\�"D��i��zD'�$G�.���&�Ox�=E�D�D�&��w��/���qs��
��K��\#�C�T�H�"o��M��A@0�4���=��nZg�F�k��H�(�3���$6�S�O�L|�2N�#���S$Ҥ=�|����C��A��'P���@��a(����E�^`����[�	� ��OH��S�MAj�2Ҭþ-���e"O�m�k�6��	���m���C""O�	P4-R�_ �I�@� �#V��a�"O�TKC$Ɗ)�$�lЋ�H�C�'[�ē�&���Y�����"���l$��=!&{�O~�"C-ɑq�� ����# �'��'P��	3̆5F6̢�Ƈ v�-�
�'�R��s��47 ���!A�Y�t�	�'R�	��U�jĴy"eḼ\y`Q
�'�4-C����%�I@+ZOx�R���Q�OԑQ�X�XzX�x�N"H�L(��z�~xEx�O���'��	Q�.���fL��%�n.�B�)���Ԥ��$�������]^ZB�	D�N��������R*"+>VB�-+ �����,=פ��F�z�,B�I'.9��!i�.$>��$�W�D�D���|J��+c�d�S@'V�B&��;ERjy���"'tR�'�ɧ�O2�9��!Z:1��!��M�
H�$��'������zTȕ q>���'� ��*�:������-es>���'	�\����Z��$���`�Ș	�'Ͳ�x� 	N�h�j��@�d�YJ>����j-�0?хHِ)�(������l1�P�s�՟L%�T�	�|�l��%��5�5�&}�� z��"U%͇[�9�5�0<1���I� [C`!}r�V�y��%#K>����0<������������	e�A$�^
"U>D��E�v���'>���S�,�>lPfJΖH�� A *J#1�(��d���T e� *����R�h�hUK�$�Ot�K���3�����y1���fT;��3P�L6p�$Yy�'
Bn�2��{���م�z\���&N>���JM5��	�v��� ��S�XBf�@dCļI��H���i՚�y��y��̟L'?9�|"�F*t��y���"�p�0A�r�������I�N�D"w۟E,�8�F�*�h�?����T�j��.Sǘ��T� z^`Ml�#r,��Iܟ������?��ڟ��	My�*X,�pI3�lݬd�$�c%�q��	�D�i�H����n]���z�#�(J��d�-�n�u�M��S�r4NC�H��b>���>I��e���q��� �����ٟ��'4,�����?�+ONE�Ti�����(ͪ�pC+�4�OJec�2(X����n���{�T�\�ٴ�?)���?�-����|��S��U��YZ�À�� �2�����	ޟD%��O��	#@>�S$aZb����R�۱�xR�rN}����6VRɺ2��p�>��'F}�%�4zaq��I�*�Йi!ʴ�?��'� x#n� ����Q盧v�\MC�'��� �(��%�I(�nG�=�Xp�J>�0�iz�'V���Ab���d�O�d�r'ĕ`D~�[C���4e����)�Obʓ�?�����D Պf���9�|
� �1�� �
O�eӁ��Rx�i#F�'�n��(�Sk�'��;m��}�Q)&H�8��H	ÓiR<�I�P�	����ʉj)T|ÐǑ�ߚ�R�by��'�OQ>�(҈(j�rU3V+�|��8ARH:�OZ(��Þ<ʠ,Zt�h��#1�?(O��8��ئq�7"ɟ�&?���v��t��$����k�(9�I����\Aq��M>�O��SNN�� RG�\ܡ�F�gʔ�9�q@CE3��S�On�:�˟�x|�0x�I�<<f���O��a��'��'�R�ӑw˄!  	�e���g�<I<�O0��9LOe�ң�:X&t�!�Iʫ0���c��0�h���pE���z��!���R�xԨ%�'�$S�������D�O �=�
p����^�pZ�e�G\���i�u��o�c�����O0�1�ȓ X��A�7J��Pb� /aG ���Q	�m��K�� 7�h�u�U4V���ȓaV-9nF?�^hX��­5�.y�'�#=E��f�MA��ӭW7X8<d�b�7���!"b�d�OԓOq�x(;4�Д@ht�I�?OJR2�"OiZ�`[5!$l����.G= ���"O �V�Bo&:M�b�:?��aZ�"OT��1��9y�H`�"��NR\�Ђ"O$�cB�0&����q�ߗ'��V�|�A �v�x��g{nm��GK.lvx��ɃH��]��R�ß���O*��cշiS
����b���ʢ"Op��"�+N���>|�4x�"O���W��/1K�08��ؓr�Բ�"O�t`�Ջ?�����l��}О�� �'�b��|�$���;p�*���M%'rў4:� �jh��2A@�Zjh<A���R�������?)�j�f-ps�[�|���2�G'�`�ȓ}�.\yǀӉ�$H��剢rD�ȓN`t3��˃X�$HKL�c�Ąȓ��	Aǀy%\=��#͕*>�LD҇;ڧq4�BReǎ�ʉЦiS�e|��.�TGx�O:"�'Q�	�[���E7u��CG�O�B�	J�4d;����%��M��B��.Fh�Z��ɂ��1�m�F	|C�I|A.�`5
W�)�^T��M�%=V"B�9�Ш�(̻�v�A쓅0+��O���|
�(�$TT)i����Bl�R$�tyRK�	`I��'�ɧ�O<�a;`�Q��ѡ!	�E58 Q�'_UC�L�(9^���R�j,a��'Y��a��;J[%$Րg�z�!�'�y��o�k�rM��"S�1 ��'�<ݹ��A<�v��pM�T�4�L>1��ɕ	e�ɗ���s3��
5����&��p���=��O�?�'c�乲���q+��p�(�'XH���&�(Y�(��Bٌ\��'�p17k���"������4����'l�x�"�/�v��ɝ�7�����2,�6����s��œ6�P��hO,�U�ӉJh��f�PfbY��.�0/$h��ޟІ�I';\�Ԛ׉݌:�e����b#�B�	�#�����OҙZ���㎑![�C�	=M8!Q�өK����ꏣQ��C�	69r̲�b�gu�9�P�Z�-D�?1�퓟.҈A�Ĳ-�#�F��Tj��R���Sȟ���L~2�����Hdm��c����ǋ�yR�!$�}JE�b@z�8s��
�y2�\�犔�$��T[$t�����y�$A��4���W8S��(�M֊�y��E<D�0���K�R��HZ����$�P��(��`{�b͠E�����+u�`hbX���H��T��e�)�Ӈ���E(M� x����-5��B�)� ����Z��٘%�ӗUE��@�"O�,���RA��(z�R%lȶ��
�'R)"U�ڣk�q�ㆁczd��'g`a'�'7[�����
:a��cH>!�I�0$p�I ���gQ=g����f����D8�D�O �?�'Q�͓ǁ�B�`�2n�,_`$:�'e�͸pA���i@R�+U���'mh�Ph�"y�ѣ�)�Q�d�A	�'�P���(V<�F��Di�h�yP��#c��tiĜ9!+�@���U#�hO�1��1�@�wa0B����eK�Q�d$�	��@��	��D4pT# ��8�n� v�NB�	)c�U3G=��l���R���C��%@�Z��bԱk��|q�L���C�I�K���1'K�51R�S��3���?����(��L�1J�
Z2(a��	�Z�l��a\������	n~����<��08S�I�X�)�A��y��ޒ"��]Q��T!C�jX@���?�y�b��`��C�?ʼ(����yR��X8�+�(2]��!�'�y�&�	�\	��E�+'�1�d����Gz��IC�B'�����d`�ɐ�ς*��ɴ�n��IҟT'��>Iڠ�X6}��y�s�J*u(p��o5D�d�$fȀ'$��ɒpj@��/.D��K�kL�p���`�D�2�L�j$a'D�x�p
�	z�����#]|�h*��$D����}�yq�������7�$�u�'�����'���kWJ��,\�3��[�3���������?���L��as˝��t����K�=��j%"/D��fJ׀M�<M��Ŋ����#�A9D�D����+GX��s��
 :��;D������x���f�H�L.8Fl4�O�p�I���(���;wfN<fE�3d}0�=9#[�O~0iC�o�t�"=	 h�'y�!�a�'���'�D��囸ru�]BR`�:4����'+<К�+\�8�K�d�,ƀd"�'H�li��6T~���A(]��Dj�'*�8[4��NCؙk�i�7������[�O<*��G��/��`ц%[9i�����J�Ex�O^��'�I��Q$�������ƛ"u�B�I���|��iA�{"f�ae�a�pC�I�Tl@yB�ξ>�LɠqFJ+H�ZC䉯K�ح+2�!#H�	���.�(C�ɋSL�s��^c1ީ��E��{|V˓����|��䞝;�������<Iz"�PyRĿ=�"�'Pɧ�O8���CJ�B$);����Ī K�'�z<��	U���vX!��z�' �Q�/T<W:F`L�}p�+�'�H��# (]H�gG�t~\��	�'Ѯ�!�����kQI�s�dD�L>���I4���I�x��{&��b#z�������8���O�?�'�|������<X�TER�Xl8���'���� �1���bcTH��' a��BN�g�q�#g�o�,���'�����E#j���j�U��T$���Cu�)KP���T- H�C%���hO`�1��S(JO>��0���|���E�x��	�����=q���q��;!�*��Cī+�lB��>Y�Eoۉ��� �F��&C�	�v�������
�,���C�	(P~��2`P��d�8&�ޢ?���%�^Tc�
��R�-�ri�<N����W��S⟬��D~�`��nB��d��te�$`���O�<�bP%_NP��F�Dg�gK�l�<� t��v�ӖE��-.�4Qh�"Ot+v�u8 ���T�� q�v"O&��Bo�=_>NI�gE�;5n0�%P�Ê��8LpY�N۲B8,�-n.˓4������?9L>�},T4���K�j=��JXb�<���/+p�ei����c-:�a"O4�����8������$!�"O�гqc��V�`��`ſ|��%@"OڥՂ�T����J^/V�`l:3�|b�!���`�(�|Z��G��@��b�0/+Da��c�����OU1ʀ?�� {��U�JiKV"O<D���.	n^EC���S���K�"O,�K7���w��dr���?��H�v"O����o*�\���V�E�2�i��'.�d�9�]Q���B��hYbhuDў�btH8�'^�Xj� i��4@�,�:�)���?��2��#Ť�7H���te�"�)����r�b�餸�6�M�K�r}��L�3ƙ7W�ɀWDVt��I��P�F�;4G���� ����DLF2/�' v�eaB�
�{�)��#¬u�����YT#<ͧ�?Q����W>;�H@hp���Y&���$_�O�!�ę�?�`H��꓄����ʯ&�!� �28�a��p��T�6��<�!�dG�@JT�`&R1ki���OU�!����B�!f��=���т�%��I�HOQ>%��̆1��0��Tr�*A�<�7-��?y���Sܧ�8�@��R�BY���b@J�� �ȓ'��7�A�LK$d�
W�I����ȓS9RAߍ��8d+��k.ͅ�B̞�I0��*��K���z��e�ȓ��R���/5�t�P���~�`�'�(���d� ��$Q!iF�j��!�ޥ� j �)�ґ|2�'���gG�Ȳ�aD=x�8P��c�sm���0Ԙ�I�>E�py���U6IS���ȓ ��8�p_HEP7aϗv�F<��2�(�g�7@Y�@�]�8>�I��I��?�1�^�':�,�%Ƣ<��!q��d�'m�qY���6%���3d�ׅ>2MRE�.7���O^��D
=|��H�V�\E $D�Xi!�ܬe�:T�CK�h^�!�F0O7!�d�|ip	�R�V�ew�)�d�a�!򤁬m�"�k'��+��T�F�$џLp��鍚�X pul��
y��g��V�bcڽ�O���O2��$?�Ş0&��pDr	ڬ�N@�<!�䆖#��X�fƕ�*��`0�Gb�<�C�=��Jq"�-
�!N�s�<Y��p��19�)ӥd��`�3��g�<Q+ۃ4�5�D��i�@�`y"k1�S�O�¸�@�A.P3L�rW�<���(O�0���O2�$!��i݂P��܁�A�"? �a�F@"!�D@�R��ѩF͖�x3�`C�(!�[,�N�i�iB�~B�����	c!�	�9A"er��F�n��Q�.�LC!�"b�k����'.V@���Y��'Ѩ#?r*]S?�1ȷY�$QG�0Ҕ�APg�ş<'����]�g��N)<d�������J���G���!�ɒjN�1ˋ�h�$�:C��Tc!�'XPf�K��ѡ�� "�!�D�)`5F8;�(�K����W��4s�¨�O@�AϜ�Wf�h�(��2�r�a��	)y�#~��Hքv4(:0h
(�B<�%���?����0?!�ŏ�SU�y0E\I#Н�!.Xn�<	��˫9�
y�穔�>�Y:�Se�<� � ���]Y޸�u�Ǳm��t�c"O��$�Ρ	��K���xr�!��I��h�z�;r>�jD	4Å34B��p�' u��4�x�d�OH�$��]��@98���`� n��%��8��( i۩v�H��Ȇ&b�@q�ȓ�h�#k݁}���C����KE�#Y0Gb����R�h|؇�6�~���_ ���ALX#78��'��#=E��EY��-��ąZT�|{b�:��؋m�h���O��Oq�&��CG�H-d�pT�&;�ka"Om0&$m���&	h��"Oت����r�0,+���) ��m�`"O"u�&��}Y���1�,�U"O�)��*+���#���X�|"� ��������E� ş\9,	S V�:����Ip�	�t��O,����	��0�S)R�@yc"O\���!6VO.�k�/M���l�&"O R�Ǉ(M`%�O7����"O���c.L�F�x��]1�E
��Y��`:��
c���� ��~�(��#�T�U0E{2K������r�d�G�`郧� �[�ސ���Ov�4�O4쨵H�	 �l����"��Q"Ov!��G8;��5��]�-��;�"O���	!m��yL٩m/ �f"OX��F�MM�5S��CJ/���ɥ�h�������+C�Ҍ�J��> juA�'�pAɋ�4�R�$�O`�.4���AN�4q��m�-�m��:��`�.�]D6��f �1�ȓLr*�c�¥1��0E�Yv� 	�ȓ $)���X����%�=�|���}�Z��B�U�>���C��FE�4��'r#=E��FϿ�JțC��"�N�@����m�r�>�f������b�x��"5?�C�O�QҐeYt��b��CS�̻���?A��Wd&TQ��Tr��
�G�!3��O\��80J�y��9��D�b
�����"n�1���_5c�^�ڡ��|R��DG��yQ�M$�&d!bB~�'�r����?���hٷzZ^�8�R�uي���b����<�ODE!�d�>\�)r��F5@q���'ʾʓS�=����#wA���U#I�/�Z�'�~E��'0�9O������Me���h	��ǘNmF�d߰+-e�sk	ز�G����"~2P�2"���`�C J�����<���F�az���BQ$�$	��i¼0	H̛S*L�=�D�W�@�d�9��'&�)��"?���Ia`��7�\��J����C�<��j Պ���A���$��!��Nў�[���J�J>��+6�]'ʘ�bo>�<�Q��Ob�M�'��o�?}�	����'`"�^5N��Rs@��=*�w�ѩ.2 ��pB���GJ��0�;D�*Fx"��F�ͱf���F���ʈ(-g�A#GN~�J�&Nٺ���Y�?#<鰃�w<�=��m�6'@`K��z~Eۊ�?���?��8�]:��i�!�4푷(���5"O�kD��r�r�;��S����'�'+&#=ͧ�?a�y'��z�����N������?QP�4�?����S�O��$`q�D�A�<�i��B�|�^��'��1ySGZ<I@6��wbr�R��
�'g$%�b��V*���*Q�cr5��'�"`�*B�`eSfM�3k���'$�����3ID�Ab�#XR�́+OڴG~r����	!5����!._�lيR�X�3F$�On���O��)a2VX�%�Ä/� ���逞T!��p��#@8F�4��0����!�d�Zú=*�+�5O	�@u�ѪR�!������{�U�u�2�xCb�/g�}���<	�%A/f�l��R#�$z���Q���T�Eun�Dx�OS�m����0��
�J�X�Cǐ�RO�麧#T�]�>Yq��5|_8U��"O���efӴks��dfG  E<jE"O� ���J~Ѳ��g�ƚ5�U�"O��!��.k���p�iXU/��Ҥ�I9��~���UZrM�u�׺{�ԝ��X��O$�	�Ot��<�$H96aq��L%Kxv @r�T�U� B�s���q��-%A6�A���c�0C䉍yc��xRV�<�"�� ��~�@B��"M�n�`�C�)��E	 fH4:H<B䉙V�\�+ŇUG"`��G3s�V�Dj����괣��N,&Yxy��J.!x��8�m�O9�e��O4�$8��=E(Y�	��!�%��DW&}o�C�(L�� � Y�K��c�E��C䉘5��zv��p�ĉ��Q"��ȓ�@K� ]�hH<�pee�3j���s2�	�6	ޒP ���`L-�l�'��b�8�"}��3�$���x�8D�d�'�̨�Iۯ�䓂?���@2��t+�h��|�C���)x�:â�?jQ
|SP(�D�'?"�J���\�OĨ\0�	�Lt��J稝'e��(������5r�'��Oe���G�x�(�GNO�!��3F�'s���:�Xf��S�:����3L�!��I"���@�I�.=P!Aڪ�k���;&��	ğ4��ןp���Ot��c*�B @T �-�D]��'����)�t��OZ�bX"��*n��O6m$��-��O�$A%�݋�~x��Ym�ޑ�O6���i��m�O�s�:���{��̒%�J�|	��y�j1T'<��'�2�'p��L���I|bt�_j�Q�b��0�ցD���'����[��y�� q -��HȽ�e�=gjr�M���I��1��5}�.�~J�@\�[	��i��
z���׬�D��`#}/�蟪A������PM2^�4+`"�O&aXq�>)��>y�@�K�$�Ʀ9Xe!�*Az"%Þbx��"T��<���Ik���|�O/&��CM�6hE"e!���AA����I@�-}*��䔆O�ɟ Y�@*f�Je�ܡ!�g�Fh�%�dyR'������H��D���E8_Q�8��V7|\(��'@(��~�����9O�l07�Oy2C�ݐ~�Bm�D��,d,��F�'�Q��	yv��p��>(�,�f <])�C�	%̸5)�y����T��X�7��O��?��X?���i�"V�Ю$��8���2@�<��Ox�O�=�O@L	����j���0Ǫ��R�Ju�
�'ޮM ��;iT`b�@Oӂ ��'�Z,9�'��;x\cD-�A�A�'��š"��M	sd�P��xy�'��Q�a$=�ؒ_�B���#�'}�� m��`d��q�^5&�8���'��ث��>tx�a%��$�m��'J�H�˞�qRM���?Y�2�';�X���(��I��^:��%��'#lr��X&�@h@S+�+\�C�'��PHk�ppsbK�,)u�(����O����On���OT�i�Е8欅�0�._,	&�Yߦ5������	Ο�����0�I柌����\���J�ztp)8q�Լh$`�J	�M���?���?����?����?����?!W�	�Q���/V�KGzL8�G�p���'Z�'�B�'���'���'j2��*gJ�@��$Si�#AL��6-�O����O*�d�Ox�d�O����OZ�d��`��e��m�?u���BC_P��=mZ��x�I՟�������I�� �	����ɺ,W ��m��"�
}k�oS�����4�?����?����?A��?���?)�zb����ϒ�Jj�͚���TD��0�i�"�'gb�'��'���'���'��U���K�H������ĐGB�t�w.}����O���O8�$�O����Ox�$�O<q2�
.	aZ`���¹"�up�ˀ��u�	ʟD�I�t�	П��	ßx�	Ɵ��ѓQ�uJ�*Ҋr�Ȥs��[��M#��?a��?����?9���?�ڦ����Vj!�Ř�:N,S���@�X�0�4�?��?q���?���?����?��(���Q�4d&\d��,NY ��i1��'���'���'���'���'Kj��j�vl�U�;E��
��|�0��?�*O:"~j�oT�>r�k��[�F>�8b	!����<����O	�6�v�$
Ꮫu%$Ue��x~�lCR�O8��p�@�'��O`LH��i�F3$�$�a3T�>��%Ö��O��:OB��	2lhў���<��%M,v-Q0�*L݄���͞���'��'�>b?9��o�? ��0l�~}�R�EL��%�D�m}��'�2Oj˧64��B��+ �`E:e�չn�(��'����Y��q�O�	_��?�Nu�X�S��8���H���*�#䋥<i.O��%�g?)�[_�Z}�h�I yZtk���<	�O2�Xt������ g�b�`D�Ţ\�tjZ��L�O���O��$��u�<7�0?�O���ix�٩��;AW��p�L!k�� ���.ړ�?�*O�c>yRj�%:=3�"�mI����<a_�(�'�"��_&a��9�˚L��Miu�Π/0�!�'�2�'`�D1ҧQO�xvO�@�6�[Q��Q��*��Y�&��'�$��H��|RT� � 
�0u�^�A%ˌi���%f�h��i�OL�$��S���@�)��pЌ��V�ı6l����ʦ��?��S�����ϓ�T� d�4*ۦѐw��f�NHQ@����'��;�lA�?)�����=��xJ�f	�g�{&)fU��f'����џ���ן���ӟ4E�t%K^pC�c��Y��LI�%ަ�?����?$Y����䟼b�4��'4՘���5�)�,r�9M>���?y��O�5Z�4���UZ58Q�3"�A��I���j�CS�:��'��'��)泟P��FK���Pap��Q����1�I����O��d�O��'$܈cJ7V���2a�6R��'�z��?9����S�	�3�x��4�סH��P��>L��0�H�x5"SX����'|r�c�	'{vl�JĪܬw|��Ԯž��$�	�� �	�����L�Scy2 �O�1� #-H4 ��|�"����'WB�'�J65�	3����OnԊ� _�x@NL�1L=���HaI�O��ą��7M!?�W*�Rd�y���	�d��y���S�_�=��(���?i.Op�$�O\��O8���Ov�4j�إ�޼-�`��TCF�6J0 ��O����O��d7���OT�mZ�<��1�HIЅ�u��Xu�[�p��V�It��'Izpl�J?i�`U�lp
C@� H�1Ӣ
��р��%0 �JQs��dy�O�"������M�z�b=`0 \�i���'["�'P��'��$�O����OP��B
�M�֩�L��=3@P�J)�ə���O�D ���o�^�&gC���"	HY֐�e,d��6nܾaEp����M�����4OZ�s���b��l�l�`��@%�?���?	���?���g�0`f!�/Jr��ALYb�g�O~��'�r�'G:6'�	�?�v%���1�B΋�Uzvy�qaӟ��	�����b@��lu~rk�]�fP�O~��Ǧ͍,rz�4
��1`���I>�,Oz���O��D�O��D�O�)�2!o�F�D�;i��H$��<��Y�\�I���II���s���Grf,Z��V1�Έ1W��%��d�Oz�,���G� զ��1�RD�A��4#���0t�n�0u�'d� dd�`?�N>*O���`R���@���! ���B��O|���O����O����<��[���ɣ������_?5����x�����+�M��n�>���?��'-��N��e�f�34�Ctl	���M�Obp����B���:�ν�p��=)ι��Ǟ\/T����'���'\��'n"�'>��3�)LG�i�GlK'oB��1��O����O܈�'��'��7M-�ɼB���Q�ǰ!�"\`ɑ*MT�O���OP�d�5j�F6�%?I1�-f���%�M�=iX
�eT�k��
O���%��'s��'���'�I���H���j�ņW���'�b_�|��Of���O���<:d��?���$�
[n���n�Ky�"�>9��?)K>����A@S�lS�E"$�ey���5�~ ZH���M�T���S�@��$)��O�-#�ũg-��6@��ӣ	�	�2�D�O����Oz�D0�i�<���'/�u�d"!,�a˄c��\�S��?Q��V)�f�|�'�p��?�v��k IR�	W�0Xi��?���&$��޴����h���O%��5��mk�$����YK4�!x�����O���O��$�O���#��P�IC�d(�B��P80H������O���O����d�Ŧm����I�	ݽb��q�P��e�������'�%?����ئQ��L�y�N#p!�-;d
©=������'n�p
W�O\�O2˓�?I��%��ԁ��:P�,�z�n�'�����?����?�)O*�'���'0o��1a3��!	�4�J���u�Op��'t2�'��'�b�f�3]Ϫ��'?��X�_�4�&J�7�8z��_}�0�?!�(ҽa��Ӂv��jC��O��D�O���Ol�}��'ٮl��@(P����о<	d��F6�����	�Ms���O������24M��;����d�'���'"��hR�f��� �m��(B�)ױi��4 ��![�� q��6s9��O���?Y��?����?)����B�s��5��H� ��h�-O���'B�'�B��d�'���A��j�a+�n(D]�Y��J�>Q���?�J>�|B�l��:$���K@i�@�� @(��Db�w~�N�0N�@�I�o��'O�6B⎔���O=�ڸ��)�-qM�M�IƟp��џ���ޟ4�'vZꓼ?q
� �(�1㓟P��%�����t�
�0��'7�=�	�����O�Dl�����LW�9��;8���� 9��6M4?y0��X���|ڝwrlQ��,[�HU ��G�. ^���?1���?���?�����i��M�t�r��=��6��O(���O���'�r�'�V6�>��58�����������<�^�O����OZ��Q J;T6�(?�;*�IՐa�DURgKT"f���c����?Ifj5�$�<Q��?)���?�W��<zE�`$�ޙB�*IbWT$�?q����~}��'���'���*�I1TJ֝��<�҇Z
Fxʓzf�	����b�)��J�Pr8��+0"neR�e�#A�Tr�Z�G+ld�'G�������|�ҋ(V�1C��=OA(��EYeb�' R�'���V��I�y�x�Qa��(��i +	)|�b|��ܟ��	�M3�r��>���y��$�cF0u(t�1#� �����?�cKێ�M��O����\���O���k�C�4/G�����oh�hZ���D�O��D�O����O���3*�
�1/V�1p���-�a���%����Ol���O\��h�dDצ���B���y\��`�,j��[������J�f�S�?rPoZy?������TQA䃁?W<Fl�(^۟�x!I�D=�D;�d�<ͧ�?�cm̱"K�q���3WȾ�[�bل�?y��?!����]}�'��'��0@��H����[u���Dp}B�'��O�YCW��<]���-�q�Ha��k�<�Z[��k��jL֓�
�C��hL�牞IhZ 0%ߚ2���bP(}Ԫ�D�O��d�O$�d?�'�y�g1(b�9
�%K���?�!S�����0Z۴��'��TCAr����Q%�#B-�xs�U:o�B�'���'���%�i�i�3���?-!ǣȺ]Av��6g�-%8l�œ)��' �	����Iʟp���������IkuC��h��O'��X�'�d��?����?yM~ΓJ���.J�?�d�9���,'X�|��џP$�b>E@��C2�Y@�ˌ�� ��N�E3��^y���98��i)�K>)(O�S��: d�8�D�L=��zӬ�Ob�$�O����Ov�D�<��R���ɺ4$��EH��w�lT;�Cr9���ɂ�Mӊ�ķ>����?ٝ'� �@���� "`��e�։��c�B��M[�O@شN�(�����T:��x��F�CV~ܹ����|�H<���'��'��'�B�'>!��ě�4`�w,Πsq%`%��O��D�O���'�剓�M�yr�H�)� �ٽ
�V4�������?�+ONA�hp��k��4y���"���Z���m�V����\>@��.����d�O��$�OJ�DN*)�H��m�V>>���� 2�����O\˓t���Ɵ���ğt�O��0˕CCq�xM@�]�w�q.OJ��'���'�ɧ��1@�& a�*C�ĘPt���s��Y�+�\7�Zy��O��L����l�	�t�6j�Bj`�r�:H��?9���?�����'��D����17���g�^�6t�,*G�O��d�O~�nY�|�����K�EC�1#Ƨ�b�����e����ɮ���l�`~��fÊ���n�<s� ���̃?8�q ������<���?A��?����?�Ο̝���DY��P��Q�1֘���/�>���?�����<�Եi����}��jg-�t.����x���'��'f�OF����i����D�_�{[�����Į1H�I��P��I�	/~��'����H�I60�p.�*д�bL�����Iן����ؕ'lB��?����?����
	���kC3@�Ĕ�)X����?9X�H�I��$&�H�2��LVz͐��û�:u �iUyC	j��X$W\�Oz���&WU�z����O�m�@ѹpaƏ(�X`a���?	��?Y���h�"�	�0p����I���6��	d�~��e}r�'�B'b����S�ai�m�PJ�tH�˂�%	\���Ɵ�����Ȼ�fǦI�'��y�i�?���}�d{�%�B��j�`�*m±'��'���'�"�'�b�'���:��,?h:A���ł:��BE]�d�O>��O`��-�)�O� ��l��Fgֽ�4͒�e�*�DfBf}��'ҙ|���ı|2P�tBۅxg`9�H�8"*4-*q"�7��$� kDFlz�jbL�OJʓo TX�*��TU:�M�
�t����?����?y��?�(Oș�'.�T D(<M:��h�R��S-2�q��⟐�O0���O�	�\ ���NG>Et!݋|��MY��fӞ�u/R���P�>�ϻ]$I���(I�)���0΀}�����I럈�	����Ia�O��QHE�]3S����"ԆI�0P���?Y�B�	����I��MC�y�JB�S�,�2&��d��гfē����?����?��Ӡ�M��O�I�Y��  �F�z��<K���"1i��:���OpL�O>!,O��D�OZ���O�%��@T�B�7�VX��b��$�O�˓O[�I�	ȟ��Oߔ�cs��7�:��d�L
��	/OR@�'9��~z��R'f��1��	i�д��⓽'�.uscIC+&��'����䟸�P�|r�ͅ%��=)��P�іa�॒6+��'_2�'���$X�(��S�? ��B�'eB83��_�&��"�'y2�'1|6-?�����D�O�I��E�W%���-�.D����A�O����<C�p7m ?!#�_	h;��I0����FYQE�H � ���a�BX������������	ڟ|�O���Y��G�U�x�b�B�j���EX���'������'�.7mp���G̓(��ڶ�S���	@+�O�+�$-�	J4��7-�>q'Ǚ*<E��S�8>L92��Ot�y``Ѵ�?���5�D�<q���?YS̅�q#�0آe�>j�N|�'�ř�?���?	�����G}"�'��'����'+lG�ݻ�ޮvz�<�����V}"�''��|"�F{���`��-��q�$�U��ɍc�VB^ΦU���(�I?	�'���r��	�����d��G��%����?����?���h�\�	N^�H���o����[	#H����A}��'�"'m�<�O�I�<�d��-����dX;6�T\����O����O����(�87m*?�;�|T���N����f��Z�� ��35V��B
9�d�<I��?���?)��?)$ե1�yC�h�v��4gQ	��$l}�Y���	s� ���7^dQIaiT-er�e�W�����O���1��IZ�3܊��	��`������	c�����O.Km�I�"iP�'���%�l�'x�y���^��P+X.O�@I�S�'���'�r�'eZ���O��D�W�]�ѩU�|
�Xjw�W�>)��$�Ѧ��?�vU���	��p͓y2�MQ�D�4��XXr����O�
��6�<?Q���b�|��w�~�;�g�YFP�7�Z,9������?1��?��?�����t쨠�	_��,�M]he4	R�'���'���?I�yr��D�+i6��H(�0����B�|�'^B�'>��q�i��Ia��Y�PH����)�D�HJB�jʘ���_P�IIy�O�r�'>�CM�
`�@�f�O#Pa�d^�	�'P�I����O���O��7��*B��e>��J�"^�f4�'!���?i�J?���hN��Z9���;D��q�С�/b�~�����r��������O���K>��	nd���#����
�*��ҏ�?a���?���?�I~�*O��	q͔�{�n��)��}����4mR���O0��æ��?��Q�������䂑���-z���V/t�d�����9$�Bئ�u7���,���Vm����* �B5�#BǥN�\�U�N��?)*O�D�O*���Ox�$�O��'v���ȅ�_Q�1�V�HϜP��O|���Ob��=���OnZ�<	fK�E�t0i���",�t��ǟ���S��w�+\�o�t?�/m I��@֑N���a������bpЀY�\�Ay�'�rnL3"
���³F��1�C����'���'f���d�O��d�O$��ՄL�J%�c���)w�}륍(�	!����O���?���r�.��cHF���}[�N]�S1Z����Gh�6	Z+I~Jg��ONc�'`e#�\ ��`���0[4PS���?����?A���h��I����`�Jz
� 1BJK�(����N}��'Yr�bӐ㟀����,�hV>Q�L�d�i����ҟ��Iğl��-�Цi�u7a�h ���͐2��Pl%.ր���U�T���'���'���'���'+��'�t��.�q��sg��i��\��^���O��D�O���6�i�OP� 
�m�xpy6�9T�e�cAHU}��'��|����/_�V	�'nD�hG����u��d����	�(� j�AƓO��q���ɥ➍ixB����E�M�͹��?���?!���?a-O6��'��J�&?jLr�L0�J���b]�J�b�f��⟄1�OD��5?�+S�q�~ة�닡q)�� �I@�@M��m�r~���*�|����~�O��.DOI��tlO�sxz��1�=z���'���'b�'`�<-���k�MY;"�\z�ȱk����O��$j}�V>5��4��'�Ƽ�'C�V�v�rQO��ˆ� M>q���?a�1���P�4���U�&/�=1Qiϙ}�uȶ
Y�
�@�vi���~r�|bZ����0�	���2�B>A�Є�J0:t8c%�^��	yy�o�>9���?a����	�r���Z���!�,���3�'1���?�����S��7i�0���nĘ}�IVđ2|a*�V��F�QVW����A(2F_�I�:7�I�Q�DŶ�������	ٟ ��Ο �	W�Fy�F�O��k��+;��Q�㝒t8�2S�'�R�'v�7-&�I�����OP��P��3c|I�AhE'=Z�%x���Ot��-��6�5?����U�n�	.���E���Y���[F�)���7@a^���Ο��	��H��ܟ\�O*>XÂ���~��E��}�BMSQ�������IT�����4�y�v�+R��9�,����	��?i���䓥�'4qd��޴�~2��" �y��#E�`ɹs�
 �?)��W����]�	ky�O!"��<X�5S�M�*]s�x�s�ˑTSr�'���'c����O���O�B��� �&�c���2EV���-�	�����O������[ Ad��E䅂:�$ZVF�qyr�����pj"n���O��d�I����z����0��D6���)�R�'*��'�2��<� ��05�0�֌�`��G�|�"��'����?i��x��&����$i�U#�8<Y�H�(�6Qzeb�O����O\�$_.w �6�%?a%��G�T��fݥ�#l�T��q���p|@�!���<I��?��?���?)D694���0\lάː����D�a}��'K��'8�O@�$Ҫ���pă��0UB5;#IDW ��?����Ş���j�#)A�(�'�P<f4(��!����*Ol�� �4�?�g*�$�<�B��/}�t}r�
�UC���+.�?����?����?����_}��'ż|;��&Pb��qGL0\븝J��'�R6�!��5����OV��f�+���.��<ڇA�x	�wEK���6M(?�%ڕe�|�w��KWԈ�UE��f�]a���?��?��?�����X�THX%Y���'�E��,��W�T������O��ߦ!�<y3#�.G�9�=
Cvmt�
[�	՟��	ٟ�"+Ӧ5�'e�HG�M�h��A�˟�Q�I� 
�)Z���It��'^�i>��������5>F���J[q���A��%D�Y�	����'��꓁�$�O��w6 YqY'^,��,B����'�f��?����S����d�R��F���}J1+���Iօ7|4 x��O��)J�?�$5�D�NL=��'�YB�ъR$;�`���O��$�OR�>�)�<	�'�l1�4n�?#l�tC؃D��[���?���k&����M}��'?,c'�J�S�Y��Z�%Ar^��s��˦�'#�,85n��?I��?Qk���v4�Q�	#���ց�O�˓�?i��?���?1������9����W`�uMP�sC�*>Tf����OΒ����֦��&8^���	�{�P�0&��]2X��	ğ�&�%?�$kJ�e�}Ă8�#��u��9�G �!#k�%��#=ܞ)P��O�O��|��l��a�!�[�6s��A��阄:���?���?�+O���'jb�'*��ͮ(h�-HKS]j�IA�@	��O���'��'h�'h�@�+�1!�@c�d���^�8@���^�n@
��x��_�b�R�<�%�O�D�>�Pq��>$ D�� V]�<Y�gD�A]�Ѐ��u��Q�� ޟ��O����OdhnX����hO�{��MH҄E%�4م͛��?����?�������4����j4y�-�����bK��ԩ�&M�N���8eH�����d�O6���O
�d�O��d�6H|�D�;��y�qӏ}{ ʓ ����L�	ʟ�%?I�ɘB1@��焄M`���埆v�l��O����O$�O1��%c�"�.�6xIu��q���&���.{�b��$�%N�{Y�ňF��Jy��܅ļ�ɕ���I7 d�U&BVi��'?��'#"�'��I�����O�"�� b-�Q�7_�ji)�J�O�Ln�B��������'-�pf�7u��Q�(�)'�������MS�O�x�#���2�M<��d�����Q���sgӽ�ht�aM�O���O���O��d�OZ#|jV)�0.0���
A���X��W֟ �I��4©O�ʓT �F�D4,&��F R��l@�%?��'BX�l����ۦE�'���B!�X�8�kPlV#P�P12��"u�f��ɻ��'��I�\�	��l�ɾ��1@#]!%Ƹ�SW�U�T�8�	ן\�'�,�����OB�l�n�#�ʚ�*l�G��(:ꍖ',P��?���S����U�
���Uܲ}�����LYU�O�|8����O�I��?��;�$��b(��׆m�T��V0:�����O^�D�O�d.�I�<��'-L;��7r�F|Y%��+z%���?9��s���D}�'C�mۃ���d5;��B�Y(���U�\�Ў���1�'I|��	�?���?I��A�%� ���$O�H��i�O���?A���?!��?����IK�WV�A��;�|(��2p���?����?9J~��C-�4O���E�V` r���%��*B�'T�|B����!ϛ�O������ J\�Q(�ۂl���'�HL�ԤXğ8�|�T������&���9�E���]r���ǟ���p�	tyR��>����?���g�ޑW�ƔL���,�	~����+�>���?�H>�jW"
��a3n�6�B��d*����͸G>�wI��=1���*��81�	�x_��0q(ǥ1����c����O����O���/ڧ�y�+]�Q,����H� ���k�En����D}��'�r@u�$� ���P�����KK�/TH-	&h�x�\��ϟ���Пxѧm�Ҧ!�'B���U� �?]��BF4!pEU*#�.$� H�<~-PT$�,�'R�'�b�'���'��(:�I�e����5��n�f��5_�в�O����O&��0���O�u��݁����U�
-�=��Fc}b�'��|���S�)�l��J�L�U���0�f�Å�i�˓0�9&��,&��'���馌J8f1VdC�d��.�;QG��'|�'���'��	����OQ�7(�,�h��ī��n��mP�*�O4EmL��n@�IߟH���<��M�p̈́8 �A��tpꐩ&KA�\}��l�m~R��<����'���y׭�9����-l,�s�H�=mr�'i"�'r2�'b"�3� �X�D*@�1��\ۄō(z���\���ɚ��d�OJ�Dڦ��<)WgF��fȂ5�À`�4�
I���4�	ȟ ���C����'"ʕ�Q�m�H��#�'�����$��,l̕��)q?�'h�i>u��՟ �I�)�$�S�T�|���IJJک�I� �'(V���d�O<�X?*p�+� ��bME� 4�'7rꓫ?i���S�)D9S�"���@�8CmD��w���+*BD3գ�!,lt���OV�)!�?7�-�DF5O4���W�XQ���Sb[�*K��D�O4��O�$8�I�<���'�2���T�WK���QOO=�Ȩ���?q��Ɨ|��'4�듻?!� �`62$�c�_e�N(bc ��?Y�Ģ�Yݴ�y2�'�l�H0��?�PDV��`o�0Z\9b�U�%�8�AV�S�h�'�'���'h�'^��{�Y`�D)Ft���*�.}dd��'"�	۟,�2��i��$Q�a<�{ ʘ�RLt��\ %U��'��'��O�>y!�i���* D:��W�NJE!$Ć�U2b�C�;�|���BK�'��ҟ��ɝZ����U:�j�Qƈ�VD��	ܟ0�Iٟ��'A���?	���?ɳƚ1V:���hE@*q�PB����'Ph��?����2vu�Q��e�`��@,�`:d{y��!wy@T8�J��4�����^f�	>��P�c�<dU��ʕ��*~�f�D�O>���OL�D&�'�ybN�Q����䒤$b⩣g톆�?�$_�,�I��9�4��'�$	I�\T�Ф�M7p�Xq�Y�H���'�2�'#.���ig�I\qVc��OF�ɴ�h�C,�(��S5��o��'������I�\��ȟ �I�<[@$X#i
]0�j󢃮}4�'J��?)���?yI~"�'�L��g��]7
�H�D�,Wix���Z�l�I�&�b>�BB&Q��zƮYo�
|��G��k`�6-N~�Ɏ
!�����(��'��I�8��CB��3&|{����Jk~l��ğ�����x���8�'ڠ��?Q"a@]�y�2a����I�գ��?Yƴi\�Ou�'�2�'p��,T����n�&�[0`�в�k�i��I�m�n�Ib�O<q��杝3���Y��/VDтG�Z���d�O����O����O�$;�'1��i�p��'̢�� H?Y�4��Ɵ0�����$�|�i�qO
L�ƨ.^Y�e�-B�#�Hl�J>�����K�7�%?�RaƤhIH`"q�� ��T	��3n�!��$�O"I>�,OD���O��$�O*�� �x?�Ѕ];�8����OB��<iT����̟��	E�dLR�*� �(c�5������d�o}��'�B�|J?a��K-d�8M�-ɖZ-��c�&��
��M�璟4�S���R�	�9I� Z����
!��q�m͏
�̴�	�����ڟ���j��Ny���O�)RV�^�7E��p&#T#.oJ �d�'6B�'~`7�,�I�����O�,a2�Q8S-��h��6y~��i��O
�d�_Ģ6m1?!q�T��~:�?��@rP���Yq�ۦ%{|Ơ�.#	���8U��{F���
5 ���2ѯ��EI�@'/oT� �b�^�W�����Î'��J�/[4�4U��	ښp#�H���̪"��c��U�C��}�v��;���2,\>�d�h6�nE�dZ��ACb�Q٢lW����H�6�����*��zm�Ě �F
{\� ܨx�}�׭k����!.n̵q��r�B�Qv�,1ڱ� DYmd���V�3�rr" V�U1��
�f�(!w"_~M�-
b'U)(	�(�!�Px;�E,��}���P">=���GWf���V'ܬ<N"uB�8j\%�6�W�*<�a�t�6Es�D�H�%*��=r-J���n���OU7��@*0)L�]�i�ǙA�lS�����{d˗�����[��3&	������J��%� <ٶ�]�??�m�0��(g(��%C��_Eh93��!����״@܉���+��2���&{/X�A��Km8�١����@u&M�55�6A��[��`U�d�����O:���Oz��'j�IşxΓ|8��i��\Qh���AN�Q6��	Q�I�4ΐ�ɯ?g��I����	۟���R�[bY>�D��f������ߟH�'��'�"�|�_�Fͻ�N�6$�2 b�Jg�J��d��6b�����L��ɟ��Ofl����
K+�e�ة7+eQ�y\��Ay��'��'n��'�ꀓW�'b��:�A_�%�� �ϰ^���yR�'���'��O���a�:��&N��PJ���S�2�'m��'\�'l��'�|$�':O�y�+�HG4EȖ�&"S�툖^$�yr�'J��'��O�����F4��9�V!�3�\�k������k�I����	�2�%�<�,�/�88�e@�?�:M{w���IΟ��Gl���	=����O����OxEhZ<$�J���G���^*w�8�d�O\�D��IŢ�ϧi���)aS(�E���ׯ$>���	 m��I�8Qڴ�?!��?	�CI�I�Pfȁsà�'�B5Bp)Y+(
U�I������iĆ��?q,��xɴ!#���R�`���h�D8
_����O�=nZ�(���������<��#�l�]2�MTN^�Y��j�+�?��<��'��ӘP*��	П4�$�[�*X�C4d@�i�( ���M�Mk���?���?�Y���'��;OL�P A:9I4`��㔪y�^HI �Ě:�D�=��d�O��d�O����Y.t�j��A@�MK��[O�O����O���'o�	͟d%�8#��?V`X��U*H�y�U�RMAyR�V&&��*���y��'�B�'T��hZ�XCk�;Jr�yb�H�k�2�d�<���?����䓡?����� ���E!\�tZ�j�*�u*�X��e�@R���y��'sb�'[�O�p�iYg�����M�'<L��2A��}n�I��0�	D�	wy�OB��U	b�����B`���͟ }�d��'��'N2���n�~�����v�n ���̖V>\L����?�N>�.O�)�O � 3�(�$�M ��CȎ�J���ܟ<�	�N{͕'K�џ�����C�%ΠR@Ras�A�H������GC�I֟ĕ'|�����d����P�	_X� )��J:>���d�
d���?����?���?)+OV�����b�d��K�5���HrG�O����<y��b����/�*E�T����W�����׊�-�Ty�'������'a�)�D��V|t����LL����&���Q�M���ӶY2>�$rUm�5hs��F`T,_��pA��'���'��'��)��O����-�6�ة9t��1=�
����գ�OD�I��t��I��`̻k�,�a�,��_8�:�a�<�v���ٟ��	iy�W>��?�S�)���#�:v@��6����E��9��S�<����?I�����I��>\:THΝu��,k�$mS��>�'e��'~�'d�I(D)��
�080Ц�q�:U��ߟ��t,??����?�����j>�"� �p�djC�ӆ���H(�O��d�O�㟨�Iwybmʎx�`��T�%z�s�nS�`o�� �y��'���'�O0맏?9�="�z��G�*s�L�x��N��?!������4���D< �D�C�60�d̂�wd��#�Pß��	ןt����Jy�X>�Iϟ4ͻBrpY���w��]�'�/��&�X��oy2�F8�O�(�*G�5��1�l��%P�ЙA�O�i��6O����ݦ����I�P�+O)�AC<+��(���K�&\����'�	����A�o�TmO��4�%	_3TlnHHd�/YA6-���'���f�.��OP�d�O��$��S>S���i�$���33G�!^�ժ���?���?J>�'L�
�̓�?��"��;9fE��$�}�L��/G�b,�6�'Q��'s��%�?���v���#S�|�� @�������'�P�	G��������П��!%�e���6��ʑۤ���E"�'k"�<�?E'�D���7<�\x!��'6�
�0V�	�@@��k���	����{�dI�t6�{���gδP����?�vW��'V�\�����\�	#�|4�b�R�� ��#��J dU��o�؀'����Iӟ��	�?�O�f���� �f	c���zc��h�d�N\���Vy�''2�')je�'�� � ��2��MI�.��L�^Lj�*нr�2�'���'Q�$\>Ь���d��G.Ābb�[޶y�E�\�<���O���?����?�"�<	�O,�cC#�?�z@8�(�@�DQ�7�'#��'v��'j�M�~����?Q���೵�ӜOa�Yis @�w(4�+O<���O��H��D�|Γ����2j�����e���YA� B7�?Q�!��<���'"2�'c⭡>QQ�	#}�F=`&BT�F�9�]oEh�d�O��� -"��|���i�*Ys�E��Ϝ�J%ȅH����i�&-�O��$�Ȧ)��� ���D�O��o�����^����y��"��^�Zϓ�?A(O��'��0Χ�?��LG��N�JF�\�_"�Y���0mțf�'���'�"b�>I.O��$f� Q���4V�+q̖BT�A��O`�O*LP�=O���<O���OL���*`,t�b��"np���WC��^�d�O\���[}BR�<�ImyR2��]
�c�* ���C�c�..`  _��y��n��Cw�_����ӟ��I�?�	�Duɕ��!>�^[�,1�I)����<i����Ob���O��SC�oV`�F�����&.�5�g<O��p���O$���O��'��	��?�h�n�b�������68%�$G�OVʓ�?�,OT��O��D�<z�dE�ZU�f�$F^L�"���l\��4O���O��|*��c��🰚���u��B�o7n��A�����oy��'���'��!Q�'���q�^�)į��L}��A�p�f���O��$�0f��D�O���O��'j�	�<q�"T�4��hׅN#FM��˟�	ן�!�&k����Ay�4��|�cb� VC`�o��d+��'�H ��'�b�h�`�d�O���O|�'�xaCD˜��F,�2h�b-���'���'u#�On���ڐwj��NO8Ja,l�q�M�� DE�O��d֦]�I��L��ȟ�تO��!\<�3��}&��bcD�j��R���뗖�P�'��S�d����̟,��8]zۃ��Z�,Q[5���M����?��?� T��'��0O��P�&��c��� �=e������$P�d��n8��OJ�D�Oڴ£Es�Bx
�O������l�O&�$�OtT�>����	,���,T%*x^�9�Jſb�u,O��z`��Ozh !>O����O��d82����Sq/��F?�����DP��}��'�'���'����O6R�pP$`ɯ\{�\��M�y�����y��'��'��O���)X��)�@ٟb2��s���C$�L�	^��H�I.3$��	-�H-���ܫq�ֈ:�ƌ�7�p=��bk��������I\���	�O�+N�"��t����.Yx��b���O"�$-���O ��B,h��=?� �d
!��5����M�؂�sW�'�2�'"Ӟ'�ö~r���?��a�Zq暺[��o@�_l�]�O>��?���)�?�M>��O�tk����w��=y򢒴uD�� ��)�����?	q�i
"�'���'وʓcw�<H1�Q5c�X�'Fj�5�S�'B�'��5�Y�MH>�*���@t�AQѪ�dm�"]�pQTǉ>
��O�!n�П<�����I��ē�?�"ǆ�A��:6��g�.�1�N��?q�Y&�?IN>�(�bT@�9O��$��Yb���:�&�ɷ�p���n���X�	ğ������?����y�@מ,�P5�Vښne�a��l�.�?�J>�a�	.�?1���<���?��Oe%�@�k���ϵ!�%[��?��f�'R�'��'�ukנ\6P{T���s!���Q��@S�ɟlCA�k�,�Iʟ �II���1Ш���ސ[�P��j��?�'�x2�'�|"�yנ6Uw���N�-;,^	sm�@�D���'�%I�'��'Kb��T!��.�Q�I+8���vgSW�� �P�,��ş�&�(��şĠ� s����HH�މ! �`�� ��*L�p�Iٟ0�I�'?)������=4��� X3m�4C��=ξ���O��O����O^l�Te�O.�2P ����2|چ�[V�^5Lژ��	ğh�Ij�������8���O,�][�zUAC&ʸ\����C;.���d�'���9�Ҩ�JԬ�U1���Q����R%E^���Oµl�џ|��蟜�I���/i"�)��A�ӓ�_�2$b��O���ȫu\���O$˓���Y�� u:���/5���S�LJ�`��rD	�OX�������I��$�	ӟ0��O�˓j������;$:���M's�I��t3z�'���E�t��$����';4����8b(�^N���6$s���d�O����Ovi�'8�I��������V��4�
�k�ꌖ'o��2q����2���ߟ�������n��-N���¤̹6�*(S���㟨��՟|p�O��?a(O�]+k�F�R#�^�a#�k����x[��.wF��r����?����?�ȟ6 ��V��n�1�AN�k�81�'l듉�$�O��?a��?�� :.�J���G�<�*PI�*���g�*-���?����?��'�����?��㎛Q9� Z��SVs�$8Q��O���?�*O����O��S,3��$Z	-�dY���<��M�����vi+�g�O\�d�O����f�'��SӼ�B��=P�`@��-!��2._ԟ\�IIy��'Pb�'#d�@�'0�<U���r��Q� �VPhŀR ���I韐��:)�����͟��	����	͟\��+%FD�u�N#9.��ԏf�x$����Oy��	��O�`s��,,H�c��(���C��=�y2�'��7��O����O��$	pyBC�2O��<i�� �
���`�g���?����=��O�T�hv��&c�������o�RZ��?�a�i���'��'�*O��$X�/k�y�V�W��	��f/y����dC�D��d�O�YK䭟pL�ㆯ͉'�"��A�����ݟ��I̟سN<a��?)�'4���A4o�i0�&⬭���.ۑ�y.�=�y�'���'Vɀ�
ɛ<*A����>ж���'���'	\OZ�d�O4�OX=�+Ȥk���S�A�^E��$��<!E��<��O�<��?����;2j�T �)��l� �P��1B�ΰ��Ay�'���'�'��4O��+u��m]�����:I��I��'�6�!!J�y��'��'\�Oش����r�"����R��Xs�2T#�IƟ��	埈�'�ɱZz��:O]��#�L^K�T�[����Q#:Of�D�O|��៞�'��Ia�D�`ޢ	T�0��]!ڸj%'�O$��"��O&�	�z��O��3S' -�Չ`��"��5���'[�'�Xѝ'��I�~���?y��2޸��!Z>8��g �4g�� �L>����?���
l���D��?��9BIh;�X�J���?�f��<��-����'�b�'�"*�<��G͙9��4; m�!bI ��
ԟ��	�ct/:�����@����feD�b�ec��ۭ'���r-�O�����-���������|�N<A�1>,�f�O,f��t�(�n3ॻ�D
L�Fxʟ���R>O.�����%��0t-Ã̚y�Mn���	���I��'��1O���)C�H1!���0������+?���*,y��O����OB�6�.6~�1�O�M��{q��O~���O������O��Ox8�R��(!J��T�
 ��D�&�G�y��+�:Ot�D�O���.��k�!
ΞR��|����W#џ��H<9��?a���Ĭ<Y0ӝqj�8Њ�m�w	�;$n̓~R&���?���?����n>�$Í
��� @_�Q)�b�O�ʓ�?�L>Q����?4��P��B������GQƠ@�m�*f���Ep 8��62]r��P�ô6lʵ�D���=1d�����i"]�'pp4�S�� %����?���?QH>)���)��6���1�T�z���g��R^!����O���+���Ol9�A��\�ۑK\�>��$ ֦O8����ɫz�D19�#XzY��aA�KU��f��y(��@W�Jb���½V���xD%UN1r�s竏	L��U8�!ifб��7m��h E�X�-�J��a� 0c��8��Iח$W���B�S`����l��A
.1�T�H<b�TQw(I6���da4GA���� @O�z��Ѧub����G (��.D,0�8=:�d:� ���Uen򭉴� Y젊��� `E�G�&,�)��A5��U�Se��:�B�SB�a
p"�+�-8Z�Y�3cH'zm���ͅUnb����qy��'��'�\p��aI�N�:�8!F� lvt����`�,�<��Sր�"5Ĳ����	�Qm4��W%���-@c}ҖjBњ�۔c�<t�$i{g�i�'����?�N|z�įa�И"/j����)D]�$:�O(�AdӦ+�8��!dR����'{�I��Ia"F���h𢈸:�L�)O
(�Q��k}��'m�Oe�i��XB�A `�P���Z��u�O$ y/̎yp�0p���g�����|�N|J� X�D�Q����h���h}��^�\X��@�T�y���/'����������V&Ñv���?���	��|��'���ڍ?�h��R�YN�Hl:����^!�$��`Ax:��e�t�뢥Ʋa�Q���I�R��Qbj��zњx�&�ƣ��D�Od��N6%G=n؟���؟��'q��N
n
��x��j�I�)z�"��OpQa aڐ]��Q'>c�<!S*�@���aë�0b�JB�a��ː�v:l�j�Dԉ>���'�r�� �򬈒oV�1���6?a!%����`������(*ϔi1Qx�~�UO��<)`��>�`YT��f^���|?���)2+O�d��ƕ�]����O�T�𼃲'�.w^�oZ۟X�I՟��'|b�'5�i] 1�*U�Pb���B�+G�>�P�6J�Xqr�Ia؞���d�c|���T6IU6�(P��omBL6$Za�ݚ�j���o��X�܀8r�^9$����e�0Y���hO�"=RC�d���q�^�^�����b�<�mI8uV�7/��o�
� S[���S}�S�`ӄb���M���?!ܴ>��P�0fB?2�>�+����[�!�Y���ɟ<�	�;���p�Ӻ%ӎ^y����яQ��5Hgj]N�'ߨD���P�.M"���6%MHg��rȑ��bv��O�c?�t�O�։z�#˵g.�)��M7D�x�ԅ��K�r����;:�p����"�OP��%�,�hQN�f���B�'&$���O.E"+�⦽����&?��	����c�*g�t���"�h�`��?!bA,�?�y*��'D~i���Q�l��a��ϛ�;F��K�O,��V�)�'P��`�U�9��M�QW��'tĨB�����H��(�"$�aI����sR��#3"O��6
ӟR2�9�F͎
���U������hTi�#Ё&�@�1@���2��՟|���$K ��M���?!����j��q#���	���cl��ںԒx��@q�}bU�'T>9!EѰR��1�#x�DjL<i��
|М�0Ǔy�$8�`ƌ�8X"&���Jљ�'���%bD�����<I���Me��t�"ճ��!3P2�r�HP�<ѡkH1b`2}ҁ`�rF��
�K?�d�)�)O0##�̂lN��I��ŧ8)h�J�a���(n��������̗'���'c���l��-��h5� !�{���ئ@M�?q�VϦ����('�@�RfZ*0^~�Q��;�O�lSc�i����C�^u&hv�ӣA�nd�f�=$� �!��0:�L��b��m���@�;D��PD̍v����ؖCp�)%F=}2�!�I�?�Hp�4�?����M[5��`v\���]�Vv�p���U#�	ٟ����̈ƀ�ğ��<�;y�<=�EՂ|�ȹ#Gd��$�ZF~��6�H�R؀�ꕵ|Y����39��T;��ɥV����!��#4�!RE?aɄ첲`�3p�B�I�ZԸ����gdN@�PĂ#����$�Q?��쑽�������q?�P���U�DM�N�z�oٟ\��s�Sٟo�?�TM��@Òlh �'ĮiED`���AM���阧�|R�G+X�Q�S�R1
�ĵ��nՁ��dڇT��"}°e�?��}��j>���B~}�oK��?a�y���V>
	 }��m�w�f��
��!�Y�j�J�r��ԕ|� � �F�<wQ��P��iK�|�@�@��;���pf��������	�)e��۴�?���?!/O�7��80�%(�N[5	ȉ��0ao�'-̬�ۓ0�\=���Â�t�T'��fOr�%���/"lO@xxe��,`D�a�H�l.(9��xBB��?
�6A�^)ƶqz���b>�Q��Ug�LC��)�0eR�,$6����A�"|�r�2� �@Y�m
%�����ǒS���+�*h�d���X��{yR�'�b7�L�!�ix�s�FXj�2}���1NJ�5��'��xo�;I�9��K��|��P����DS"05����#Le��m�	7Sب��D�	�����O��D�<�Ϙ������5�4��H�?��zQC�A�<)���&d%���H����QX�D�զ�Ioy��(m�6��O��~���@�E��D�9ф��7����Ky��'gr�'?��(VB%0��O�ʌ31�i�	�%^���"3�Ʋ>U����C�_2�-�}BE��)+�H��dˋv	�Iǉ ]�'NY���?i���?Xwe���F�>mȐ[���3ft��'�b��Ӷ9l��9���a��-	��I�)�����~?Q�ۖ*�E�2�R�{P����
5��I�f�mHݴ�?�����'�?��4h���5�N���6�ރr����&�'�fh��'�1O�3�ğ'gv�8@�١G��1Є����	�=��#<E�����1���.��@���MZ��$��tR��ӕ �\�#��L��ȆeX�p�pC�I!�(2��\�'�����!'oj�>�e��;+i�@feQ�xQ�|�n�O������?���`���d�i\��'�]�\m�:lj�Y��^�X�a��N,;)�O>\���'��@A�,5�:�*�3^Y�݃H<����F؞��U{�Bd9ch�*G�L����:�$зU�"�',�a�kA%}���H�l�Y��'](*�#�+�Z�{��0��I�'N�"=E���ڤi���R�"K�G���y��P���y�D���O��$�<q��?��O<j�R޴X���1Ȉ�\d9���O�����	��.7��*;Z\;DP N���{u���^5a��F��M[0C�v�8��'^�=�́w�Д9�|b�'>���O�*pJ¦�7}�j�@b�;\�Y
�'��$�� �F��Lx�5���	7��Ī<�C�3o���'!R�i~VMi��-+ ա���5U�^���g�<Y���?y��U�X#�Ř�u�@'b������� d���QG8��O��p0�S�#���f���p�
䙶N�=&��#?�0,�����~�fK� ���B�;<,��	Z�<y!k@)E|�4����4G׬�*�n�T��@ �'üq�$K,]>���`B[~�B
�'� �S�
XQ"��E��Y�ֵ
�')bx��Q�X����B�$R^��L�$2sgD�.G��0�Ʉ�H�r��8�	5�i�@R*,��A��Z�6�C��+�P����^,tD��d١*�TB�	���)����=����O�&U�TC䉸.2����C�P��Bĥ�y_nB䉡�dY��H�ln�t`Z62�XB�:~�Ԩr�B�f�L��f�Q
B�ɸ�Ɣ
�K�[71ѓ�%��C��-i��a� �*]k�i4cʬC䉶*�:,��ˢU\rCP�� 	nB�I%z�!����2tH!�*�ϰC�	P,F�r�G�>�t`+͉=��C�	%��6������խ�3XzC�ɬ ���S#?��)Sb���GC�I&W@IZT��5B���U��	��C�	�AQ�xk��`����cd�k_ B�0.ʵ�f"$M#��FKB�ɓ
��D؄�-|;<�Sq�F`��C��6Ψ����<�Z :�͇)T�B�ɳ:�쁷��W�՘ ��"4[�B�I,zPD���ɼT�9�J ĲB䉁u�d� Ú�S�F-+��7Z��B䉩y��(����t8�Z�S��B�	QJ���'M77"�̸6�!��B�	�\~�SAXL�ʸ��,|��B�I�>�2���
��3����E�1h�NB�I�5� Q$3)Q�!�4Vv�C�I�"ͦ���)U��Q���]�C�)� @݋��[����\"�a!�"O\����? n�`k%��yؚ�"O�,�чܒ?��H��(H�� �"Oͳ�V���'�L�}��ؘ�"O��[��ؽ��-BA��U�����"Oj�)@hθ9oZ���jU6mcn	��"Oн�%D{1��r+SLmD�ؔ"OL��ƫ�t�YuI_�m7�(rC"O���E�J��|�h6M�-���h�"O�8Q�l�t&�1#��Vv.e�!"O�]�w�y��0Z�W�Uh��C�"O�<�pFЫ	�
^�9\�U� "O�䊆N8�>}���Z?&C���"OVm@��O&,�,�k��X����"O�V��/Pt8�8�@=`���6"O��;�
78� ���ߍ;�% C"O�%bf�͘uA�������V"Oz� ���6��z�CêBli�"OĬz��?l:��C�|C���@"O�8ˤ��!��'��*}S�]�&"OdiG�"O���X4M�u��"OZ���g��'��(�vi�0R1(1��"O�E��o��<�b}3���	��Z0"O�M�����Db�f�+~U
��"O L���K�\LQ௜�?��A��"O�DteͰ/�8����/{�%��"OpƢ3%�|�-߸k��k�"O|j����/2�s�؉r���a"O�5z1����F	 bn�Eb��p6"Oj��ңV�Ј1��x�P��e"Of�q'C]�x�D��+^�@tܩ��"O��W�?S�MHS�TR�,�P"O����/�]� q��a�P"OMP�鑸m�64����3�`p�"O|-�"��!���H2�@ e��PF"O��ȅNJ���X�j�`�bS"O(TzDHn�xtã��(;��=g"O0,`d�IE��SB,�<ap}p�"OF��$ʛ�8�d󎌤C�"�K�"O`u�l[ v��c�[)q���C"Ojqs�o�?hI�=PB��Z����U"O��� �F��������aG"O�y���!B�p��"t�$�"C"O\ݐ��D% A�����^�~C�a�b"O�ݓ�ɔ9��Qy�	�/�b�c"O,���O_'	_b͘bB�
@�h-C�it����lx��$JFgD�
�ŗA;~a���6\O�a��䐏]Z��P�2h�E�[5H�\���В$�n0��L9��SH�#`�� � ��(��'�h`!�`t�4�M��Q?�`�H���9�H��m���8"�T�<��%f+2�`�74�� ��-PV�Q�bc��(�֦Y ����M?�䁡U�3Ȫ�R#��3Z�2��v�#�Ord���ύ~�ƭ��"�K �e����R�v,���H"��ڤ���z�Z�#�{R��}�'Q�4�+$G�|�V���G+@�F|����I:�D�j�4$�ȅh��ԓg1V�Ȓ!I��j�bh�o�	��`�2"(�o�����%V��0녮�1�$�w�XJŀ��
�J�Z�+ I.h����i�q���S
B1l�9�
���i�A�3:�*<��W��IR1Y��1���6{�Y(��ނ� ����U��X3�Ǻ�w`�$L�t 5}Zc��КcW�5	bH�R�Y��()�U�<��W�`�*�zE�p��i�D+X� 26+�[��W���*@P�J�3A��BܧY�JX��cM)r���վ4��E|+�O^d�i5�A�5�n��ߦ~��"�*G�������b���bC����
0�A����g��R�'���2E��#�%=JT͓%|���0��~7*i��@��(�N@AO"l�H�@g��?�&T�g�|H��qa�ɕ��?� I�Ĭ�4�xȢ@�g��C�J�^��,+�}�0�91e����쳱
���i��)rƖ,j������ߏ.�`��(�O"�s�-_��u�Q�_XA#Su�$ٕ
�X�%h�eյa�Ā0�'Q|�
�hB���{SE�V)d�0Gg�5A���0�)�7W��s�"�	qq�M3�M!zG�^r��S�˱m��=�e��g?���H[�e�7M/.<��d�:���+B"I0����U�ߌ<l�9#'�D!S��\������I[�_����� ;���6*�)�]�慔 ~03�#���Px"��%(��-i4��:!;���n�x�]���G�μ;�#��?�ه�',��!�O�2?�HK��Bm��beT�Հ��'�p�Q)�j�����!``-f/F�2:��Ш-|2T=z֦b��[�j�4,,�s�hcj���j����G�R�Ҝ	$�;�@��@����z���)G:S���,估���r��@p6cS�J
��Γzk)JK��d62���ͣc�����Y��hQ�A����a��סB�}x�4�ҠBܧ9_M!�� )5���|tΉ���m�5(�b�<�'R�"�d5b3fL3Gd��a3�#{$]*�-"5d�#�&�2.�\PBgS'!�f�'fT<��w�z]�gO.[l��%+�>�pt��YB`����K����u��"Z�L y�
T�HYi��\p�u�D�u���'���$��%���y¦�'�}�v�-N�Z�@bS��OJ`*gM�J(t�Fm�7_����7��|zu�D2_�j�P�E��
#f�`��Y?	w�3-�4\	�x
9@�)�5��ʦ�E9����ЂW���9C��jaH�������O/F��1�x��5��8`��3�'Ɋ�=c'�9�OT�������~�ɇs}&$"F!�'ku���� �vx(�B�`�Pꖇ_?f�xa�O|ў��Յۈ�2
�2}(Ō��'���H�O@��	5M@)�Q��*2@�`�,'b���5� �F�Bu���6�Zb�Hzx�Tbɖm�f0�vD�'s�r�2�$56�p�v(Fcyr���C���Z"��=i�i\����w�����H�$M�R��7�ܲ)��3�'I��qu�ބ9��@�M�h��r�d�W��y��@
�$}y�/�uWFU<~�XS0��v��Inj y#��.; �k�n��I،���$z��}��IZ�U�Re{�F�8���}b�5��mU)CQh�WK�;f��FXO�X���hO\�ã�6��!Z7�[W�ԩ����v`"ZЁN����+A��hp �+`j%G� {{��k5v�b%2��Tv���5R.�u�4�ŌO��91q��F"�Ds%�[4KtV�$�h�ƊĶk�ꬰ�i��&$��׼����CHp��"H;ܦ��qALN�<ѲOٌ+�P��B�/m���Q��П���b�X*v���GK���ٍ#�x���.��sӨĀ��ި/������2t�!�'�^�Q㢐�-= T�I�QV�eť^NPi�����). =���^+����'FnA�M�5=�|@�h�\�l���+����̒��x�)^
�)�u�S�}�X	%Y?_�Q�*R!�����'c�8�)͍H;*�Xr���y���%F��r���$��:U��v��Ĩ����wT��G�+A��8q�G6kv�d)�'������C	�`���U0n�N�Zݴ?�a�P���S���]�P��?7��y�����.�ث�N���!��9{��q����%��NBR���w�'�^p��Q#y��tU>�<at�ɪ!P,5�R�5n$`Se {x�dC%�K�D��ڧ�?м)I�-��B�q��lIU�cm��>��� %2��6��U�R�JM�'�lи��ND�a�(/��O	���u�ا[��#ՉT�vP�	�'�@��D�_d4��a�%~28<
ٴ�ݲB��^6��χD$�~nZ&z��1G� ���Ie����C�I�HT0�� K�oq���s-މ%��1�價�ލ���;������IV4�G{��Wf�+�M�$�<K'�,��<!�͆��(cW��f"���0��, �1²�[0>��ၫB�P4n��� ۢ.��}�O�9a�*y�VG�=��i�����Xyb-��V<"��aP��Y&Iۤ���W1N�d˧g����K�6���G� 0:��������v��=V��r�IH�Mw^(�1�lod���ŋ+��XД����O@"t�S`�U�E��>�"���I�e:ވ)#(:$��ˠc#
J�e��-�����u8�YYb E9TAv}áZ )�Ly�#��O�$�!c��X�=��U>ZJ�XC��'��+�I({��H�� �?l���h�v�y�A�P�P|* �	j��Ȑ��'zı)���evy;��̴�%QL<�&�ɛo�5*��97Gv���,�)r����"ۈ@$�Bc�$)��B�ɨ5�=R��^�
kH�!l�O�j�
	�"����(��~&�� C풒ȶ�h4Bב-2���F=$�T�tᅢq�8��@��V<�<9����mR4"Wo��<\��)� �<�BL� ���E�\>��d�%�'���/�<��`�'Vp@���9bv�e*�(oVڬ�'\x9���1cf��� +̨)9��C�ykL�(;��SR�Ss��uA�NT ��x(�<�4C�ɩ2�0l@�h�|@,8�!�Ǹ8 �B�	��^(;%�Qqp�����C�*s��؛���3E�:Y��hÈ$�B�	>sX���ˤ>:@=�EM�1��C�	)?cM�FC�.#Fi#�Y�YǌB䉲Eub����:����p����C�:�P�`E�Z�-X@��;s��C�	�%M�r��	d�t�q�F7r��B��F���)�`"��#��I�'�\A�S�;NB�R"a�[�X,	�'��%/Y2t�i�O�WD"�i�'h����Ʌ&��X:���@le��'�jHlɛ��x�e� ;$<��'<�9)�K���x��d�:���1�'�J�&�_�PQ$ ��.��)��Z�'H�%�T�^)Hg��B2(py�'���g(B�]��Yy��*RxZ
�'u��!��=�\�Q��V� ���`
�'�F��m��n7��Հ��Oh,) �'ƈ���^tE�p��R�x��'x�y���In�I%؉^�4Hp	�'�f`q��P��Pu�ԏ��YtR�'�R�Z7O \m��#�D	U��9P�'Y�೓J�/�=
�!Ե{�r�
�'��D�4�
/�b�1s-_���؛	�'D�x�5nU/���R%�R���'���1fhˁ!��X+%�Q@��I�'��U��GC�x��:V��2?Lxp�	�'E�@���%�ޱ*���$.���	�'8V�IC�y`9�P����'�m��!��0ìH���Ŏ�Pak�'X6��F]bQ���i]�6����'�֌�K�)>�!����
!�ꔡ�'��$c�$����	٣�G�*UNP�'���X���;G�0X�^�&ȒU�
�'s�Q�>J���#���K���
�' $1p��O�m����!
�~ZD\�I���c������A���1G�?�	�F[N�" /�#<K�����$��B��4q4l��Ċe�(�2 �K�ОB䉆+ �$��a� L�b��#�$75�B�	�l��,���O�!�ꉙk׾1P�B�3Gۤ�'���4�n�.�B�Ie�����e�4��Qb	#�B�
,���"���=Ls�x�c�F�*jC��-p~��P�g�BL�����KCC�:W�ά%���r,˔� �M��C�ɶ�x��&��$Bf��%�Z�E�vC�	�������M7�&�R��7rC�	�c(x����(2֭[�
~
B�I�FǼ�V��)hP�˵���i6�B�I�q<A��B
sK����FS�+Q�B�I!ll�l;���1�P�E��B�I�G0r��@d\�6vX4yԁX.�LB�I%:JU�7��2�"��6��8�C䉽��a�*��x� `�U�
�3S�B䉸l��-PT(��Ჴ �$Z�B�93a�q���}s��.Y�hB�	��ШpT L�Pg�+�*B�ɾ0W��6�Q>5��M���� r%�C䉖 TH��{�Y9�Â�A��C�)� nD�P͇;��LXClQ&m��I4"OV�ـ,J�rD[�ۗ����"O��wDB.D�́�M������"O&�
�m��N��١d�4�bD�"Ot@���9wj��k�"Lo_�D"O�-�F)7�\��۫Y<�)g"O��i�B�|g�4�K/=�d�"O�̐��B�6բQhE)�E"O��i�-S�p��z�9�L��2"O�5
�AJ�>�����^<8�0"OfZc_k׮�`Q��!=*y*g"O�8ۣ�
k��-B�2Y6N3g"OTe�cb�XPd��Y�=H��"O�#�j�'n��sc��{R�LH�"O����	g�LȤa>0i��"O@���M["s�����޵3�ѳg*O2���g�2���p���F9�ybǘ$T��#s �)֢��y��9U�j�k��fW�ضb���y2�R�r��(�gI�WE~�	G*˙�yR��)J��8�`�'D�*��Vl�=�y2��yn1�5*5)T�(�kL �y2�z�D��#!��!���ױ�y� 
70�a�����a��#�y�.B��,��BA�܆�sDf�-�yRJ�)!���,�<$Ӗ�Q!��g� aA�ˠ��i���'"O!��ĭt�̫��۫Dy~�*���T1!�$�P�:����#dB1��ņ;!��T�[�j<I5�P/?YјB �m!�䚻�jš\�*4�ĪŎU!���,����l^�33�!�7��?F�d�(j��"~
GN�%��#[�?��5E�C�<�c\	=��$��k����pR��{~rM�Y��{�m��K��&��*D�"p���ʯ�0?9��ֵ�?1� Y�05*ăN�]w*M`*�t�<v�*�be3��N������b��ٓr�p�}��`�m\��z��8P�ݸ��Qg�<	�_��6�rd��EA }�bk�<iPh�.����� ZDJL?7C~uۡfB�|ڥ��"O�)���.���ŀ��d�R�+���~�-�-��D�O���$��G�"�䋭`삄�D�P�QQ�~dU��?��c��[_ru 6`�Ƹz⩔o����-Gg�����A�/�T��N �9tn��Fg*\O���b���DV�*B)JF'�2&EH���ćRA!���;��1�-$��E��fA.2qO"�k�(�%�0|�� 5"��Z"5��x9^\�C�	�cۼe��C����@)�D�y��P:��+�Q>˓~Gf��2E['s%ҍ颏�	m$��ȓZ1��Z�@V�i�>��`�zl8̩k�E�dĆ��=sk�sa�O
5�؁s�nY$$`���D�6`ܸY�O,P��ǭ3��|[n_ t[��!�^��smPz�L���;u�D*$�=���p�&9�> �x9Z���C��ɕ�L� �!!i�$����X�dC�S���g
��gjn}�G^3�@�3��N�=&@8z��Ɨ��T3��9@��S�:�l0�+ �1�ʨ����ip��!��'�$h���T�0�i$��4���$������Aٴ<�t5��O6M�v?��(4EFh6H*"ԟ0`�W���F�$�V���+j
I��C�&��O�XhpB�*E:8�������m`T�'�n�`'��CX�d�ɀ)�j�B��V@�����hU62	H(�)���O��R%�� 2r}�4e]{<س��O�3���ih���Ɏ�E�z��B���L>P�A�3��k&阇Y�
�aM4A�;�d �&�x��?��5 �#E�\-r<�Ӎ@#|�����cM#��>ͻl��`�dB5�p�o�3c�d��ɠi�ƅː%�4L�"t���мF'�JQKA)6�$����48E�D��J�3 ��
�:�� ����V O!�X���|�v f�	"!����F ��Y���"<Qv˓^��+��H�/ԘQӰa�p�'ߨ0��i�o�<� ��ҵ>E<���A�`N�s�f�'.5��0lƦ{��	B��x�V�N,3@fm���1��z�b�#��˓v�HZvG��B��\�C!�ؼ=�dϘD����aH�!FԒ�/҃kgX��.N�9���IΧy7�%c*^�ke)�/>.�5��"�p>�0j�8��F�@�D�T�I��?vx.5��+ȏ^�(�E�/I'_|�����`�zР�/AU˦��@Ǖ�{ ��H!�&������X�K���Fˍ��4�K�<�$��:K5\!��oA���Q7k�
C����Or�#�fƌUv��C��Dx�,j��I�۰aCQ(U��z���ޏA�h��tE����M~��@�Fȟ`AU E�Hoz��޴��FA6�U�cfK|�¥0�ˇ�|�``+O�z�5���'�"EÔ@�4!$����W�8K� sE!B��DJ
_��%�� 2wTў�]`;JY�����ON`�1O�g�b��d�[�K`_�?/İ��U
B����e���o_����FУ<��M*���a���/�����N+{ޖQ0��)<o�,�7T�'}��Gz⮇��`��W��͘&ĳ~���񲄒 02��b&'�aۄ��'+	��A�^�����NS�<��EFx�+_" �^)��Y' 5HI�F�4�r$v䍲p�tVO��q�K�#O¦�Pʙ��j	��&��T��D�7kvx�Rվrʩ����P^��z�n��o�P��%�'CjE3��3���$a�si���3�Ns>\1�o�9iZ6xqb��jD1��4�U��-�n�ęt� 6(���T�'��(B� U�j:U�P��_�>=�V	Q+[a��!@G��m�.M����3H��O�|y�
�6��G��u[�\��'M~�v�B�%c2BH�oYQ���A`��.P��-TF�E��-]<>D\ŉ�o׃ �|��C�ؿNq�yÝ��H�@�?������x���x&F4 L����j%H<rE���0���Ʈqh��r �싂�FZ��EXbX?�ccWLv���2r̸�s�[�l��D��}#'Ϝ�~��4���'�2�9�
B��;SN�:nb�x�#۬3o �{T���S-$�pf*��7~2�;�R��h%I��?ͻ���i�.�]�ӏ�$$ ɇ�	9(2�Ix�+I�"/ܕc#A,�x0�kE �E(��U)R��"��'.J��& 6C�<�O�
�����%Kf>�cF�ӛK��Ba%PܓeIh��X-|�X1��^^�[�����i��Pnm+�	�.M���GC��d��n��"����8��Krb���*��*w.<x��B�`4����:���p�ʒ�-Y<UI�k���~�O,l˞'���@^=�y	�B����!�h��m�h�a|FM�Hf`�	��F�!��"7t�!9%�P 
k<t�'ˎ pGo
r?Y硛 ����''�Di�g}2⑁�X)B�n_����;�G���O�2g�!#��R��͞>�FDQs�e�F=0�J�9G>L�F����fpC�f�9iBD�s���*���.3R��0���S� Ep��0&O�^�PI��nL-SZ���X�aM�=򠐦�͸&�q���Q���)�O�9�Q�v�2i�!S"��*=����o%(�~!�r�'���0��u�n��,*d��ZS�.C	���G�JG
��|J�L��<9�4j���X�'����f��;h%C��Ց`��9i	�	��$۶�H	Y�L�RWo�2j�d0UjJ������ŊP?� �����5aj�,[BU�����ܬ��	�AG�%ʀ�؃M�I�P!��3�l#<���/��	��G ����R"��@5��^��Ī=3�X+��� 5g��lڐXt��k��Pwn)[ޑ�D����3�da�����Lq��S�+�c�L���Y�a�4w):D��ɋBFd`��}�I�Snl�e�Ұ\kp4���ߛ�0:��&�O�9ZLţX�
L�+�%`MڍB�ʏ�u@T�1��e12�>Ҭ�4*�-���:�&�$���Pj�3!��O�z�\HF�U�s�>�BB*S+�0|Fz��C��.%!�"ܙ�X #�������F#Rh8l�aK�>v��h`�0|��z����>���[H�{��0��[b U���2&NG�a����9��('��8F��*�./�2l՚��%�f���~o���=����wI\�e��m 4)C0��e�7"N��W�M8>޵
��@1�y!��Y��?�T���]��d��DJ�Z����&��ڨر^6]ͤ�`ؙ�(O�$�����:5haӇ�D;*�R9� U�<��!A����1Ec\��� ×�M�~�D�<%����3=&h����p�剖 G��jt-ץf��$�Ac?/�8���Ƕ$���)	����֫0X<i��U�h@��²��Ll�׉ճF}a}BJ�i� A�C� �E�s*¦��'�ND�5�r!ph�2q��(��t�T��-!�e��`�����b���y E;g6��V����]9� �^Z�I�mM:��H�"~��<��UY��!NE�s�Z�1�:C�ɀW��!K�d�0��)��C�t�O��Ӯ҅��<9�U�i�5ꃥTvҬ��ft؞� �O��M��IPU���ĕ�ԸUφ�YcD)PV�14�8H��	�^#1� �0ܲXɤ+=�	�(^"�
g ]#pj� ��� ���7�A;3��Sel�bS��"O&0[�'�]��\@!��!bI�H�k�o�� 4�u��nԜ8�fq&>�A�je�&�>r@��#�@Y�i�r���	�v�+�]��;+[M�c%)=�~%Cuo�rE� ���g�4e���m��ܪ�]�J�tqWAV\�Qf�.��Sq����x������}���A�F�<���Ȏ�F��䓧�yB��O�& ��T����̌1�,����d�Z���E�?�v��U�д7r��2��b!�ڗ2���ǆ ;Yv���t$֘A%b�Z�~d����W�)�1���-��SP�0H!�)@|8����{��}22M�_�!�d�D��t@1+�P�D���
���!�d�:���T�~��"'ƗbY!�D�0?��1�$�>�xC��P�nT!�O=��$L�v y	g�#�!���}j!cγ<a0��V�d�!�D��hf<�5 V42��(�r��>�!���lvt)#gċK��P�D,'�!�$�H� �s���1�2��!_�A�!��'��պ�l�'{ $�� [/�!�Dqa�(�T���I��ڤk�0	g"O���F^�2ݓkU!?D\""O�d#a��V����	Ҫ@�t��"O
��UL��sHF�� �î#��5;b"O��a�-�E��HQ�-�f��u"O|с�`�	xo`QIׁګ��Lw"O̕Y �*Z����ݭS��Ԙ�"OŪ�m�<ko��+��������"O iqQ)����.�:aNi�@"OD��a$[�r�J"���S�R��1"O(!�F�^�C��`,_$]��@/�!�$�^2r�{U��jW�T��D�/�!��S�{UD�0��
��PWDǁY�!�V��nT�V+� ���Ӭ�3I�!򄋾fҥAA@U&K} ���
�m�!��X�	����f�Y#"m��ꝠQ�!�DĽj$�3d�MU�p9E(Cc%!�R�eӠ�Yq.�	=t��	 !�I7%�8�*�'X�(��4:��_,\!򄅚F�\3��I��]�sbوt�!�ռq��Z�[�a�XE������!���N�X!*FR�;l%� �=1�!�d�<qˌ�x��V5[Gb`�Cf�Ui!��R�< ��aҁ��%1F��уdJ!���gI
����	z�H3�S8�!�ի65�l�	A$YCr4��ٔz�!����a�Ͼ`&�1�a!��;�!�dZ�Z�ZRcծJ�U@ k��v!��1�VTS� �\H��$z!�DR��p��',�<I�v]�1o��!�PA�,��oߜ$����IU7!�!�D�~ۂ���B�3rp�!�8�!�d[�3��<6m3Ь��I�k�!�Dd��Qss�	�q�j]��B��!�D�aD��!�@@�o��aB"_')}!�P`�L���\�H��l"v�3%�!��ݚW,�QDKP�D�~푦�ψ�!�$�_�P��Q	����]A�a�,2�!���$�~�R�O�%y��1��@�0�!����Is�F�.X�MkG��s�!�Ĕ�9�f!X��L2��Q*el!�$�<�l C�A��,�>��b 6s�!�H�@c4� ���2��|*�b��=�!�P8[�^}�a$r�J�Å h�!�� V�������1SVf�+���c"O����15���Q�4�|��C"Oن����xrT�Ɗ�jH1�"O\�����4��C�	�Z��1"O.����L�z;b�Ȃ���=S��"Or �vf�r0��� �d&`�u"O2�S�5�n�k&	E}�:(ys"O ��
P�I�:ŊVj�V��1�"O �AW����X� �Q�[&�y�7"O �bDE��+h�\xG�$��,��"O��ҠjÄB�d9���D;f�B<Z�"O��� j�{ 0�jpg��`��"O��j�KC�~����(T�zŞq�"O����Z	o�D0h�&:����$"O������B��!�L�f���"O��J���'u�Ѐj�BM�*7"O��3��\��;�Z�V�H��"O�P �0YJ8�'��`S�,yD"O<*FĚ6`�@lrk�i�\1�"O��S��d����N�z�f���"O���j�
)�fɑ�� o�F�ҳ"O@� �逑;����K����jf"O�d���â<�$+�o笉��"Ot�
��8Y�H�ywJվc��9�r"O=�A��Ek��CDL�;1ȠY$"O�!�w*W�p��Zg%��$��J�"OD�%ǍOc:�eDV�R��Q2%"O�0��;!<J'Đ�%v<���"Oƌ��T(i�
hZJL�����"O�!�)�"z�Q�c}�fq�T"O�{��;d�اa��( ��"OD=ÄBөW�U�`��^0v5P�"O*Tãc�%v��8��D�E�V�b"O`�ʂ
R\�# "S�9Q�"O4;�	�,An-�.]�La�@"Oh�z��M+O?��u�	=,��)�w"Oxe�r$� ofH�S��5&�2)5"O:�#�m�B���������58&"O����ވI�f��e�,sj`�²"O ��k����Da��Nt�dӗ"O�� W��L�� �/��.q� d"O�Z�H�"XzB�n�68x��"ONM�1O�&�b$�TNɭ�I�g"O�I#LC�xw�0�ө'�d�w"O~�(��;%f�D�'-�c����#"Or��T���.� =�Dɑ�N�4 k'"O�+cZ�wk�!��Q�f�Dۧ"O6��I��A2h��fO�yXA�c"O�h`��&Kg�p9g�S�E8�e"Ox(Z�e
A�Q#��&3�� "O����3R��J,=G#P�qp"O�"�
�][�J��Mt"0���"O�$;#�QO7 �2*V�+HD�0"O�5���,m4��q�(���r�"Oܑ5,�{���I��N*�r� 2"O�0��͊�W2 �ÀA�(���R�"Ox� %O4����3���=�(�"O��zv@i��g�3u�`bW"O��f�P�.6^Š������Q�"O��Qu˄�f:`�	��M�D�b��R"O�-Y�\�:1`9�85"OD�Is	��\da����fiF=bT"O�4K�YF^9r���ZTe��"O�P��H".\]b�a6<A�E`"O� h�#��A<�|�0��E�k�b�0"O���uI4su�H�'�N�����&"O�td	�4��DG�����"O����퓺C�Xf%I�x[��P"Ovā�y*j��E�8x�Aw"O��1�̆-/@,�՞+�����"OV�Z�3nU~h��oȵ?�@I��"O���̶Ok��nS�v��ٸ`"O�D
���:/�%ɡ�C�U1��I�"OX���R�P�Uzvo�m��)P"O
���#Ĉg��a�턌1�\��"OJ	`Q��;3m�0Il\0f��d"O�Й�F�l�N�����1�z$�b"O�ѱSl�dڀ}�%�W��8�"O<Q��.��`Z�J�W�<d��"O�mp�G�tD3��`vAb1"O�N��j�؁���'r:�;�"O�����F�]�!!д1�ꄣC"O�x��C�t�qq�oQ	1z����"Oi��h��[��n
�i0	�"O�����|��9�̎�C��:"O���k�%�	׬0��qq"O~遵lU�H�X ��%,D�$T�"O <���T�N�(a뗏Šg�LI�"Ox���!��8X�.ȍy�\8rF"O���'䕋1UP����Z�;z`G"O�y�3�<d��� �ٓN�U�"O8�ҧJ�F�pƊ�` Y��x��)���YY�� ͘B�0az㝐3�B�ɺ���P� T�XG�x��?�B�I�{�t��F�&����E(�C�ɠb`�Ն
�������ǜ��C�ɤU�$T�'���9x�1���ǻ�B�Ib�.���"ArHd�а�CB	B�	� ��t��D_�f�~	j ,#��C�	_�0�HB�3yyf9YpC]:
l�B�3��Y1�"7BlC�FI�B��;M����4(sCܚb�E�dB���  �VoG�oҺ���C�1b<B�I"i��Rf� }���"��\��C�	�T|���%�n��L�O�C�	"���k�`
�kmx��� ՚O��B�ɑ[�p ��ɿ�V�a ?)g�B�	9S*�a!IC4~di� �CHB䉙`�؝��I�S6VDEkM�A�B�ɔ1�n3"�4N(*T(�3tD�B�,X��eC(O&� �xB*�U׾C�Lq< ��Ǖt���Q$gL|C䉳�F%Qf�K����i
>�2B�	,w����O68��� ��y<
B�Ƀ(�@���W�Dy��
�+$C�	�o�N X���&� 5r�*����C�	"y��
�nũk� i1�	B8](bC��(�z\�%H�.Ŧ�"R�^�B
2C䉰1#6����%�R��e*܄�*C�	�#B<u	�#R-0\jC�yFNB�	]���8sƄ�ZH@q�dG�M�,B䉃��sfbX0�RH�䆹v�JC䉂o�2D���
u<��W��r�>C�	�vj7�Y�.P�@�BV.�6C�ɻPŮEx4H)I- T�!�,&$C�";�$���/S��p
�F�B�ɕ5�Rٲ2
�J��ac,E7G�B��:����B!�Y�:U�v���`�:B�)� 
la�d��J�T�r��_���"O�%��ȅQ�
DѢ�ʚR���"O�i�%��؝:���)�3F"O��h��;g����P�7.��T"O��HٳJ��xxag��E��A��"O�P��96�UY��[�N���"O���I�}Ю1+�@X�R�ν�c"Oh������t�4dat���2lp��"O1B�	�!{~���IՐ��[ "OTP 嬟""�PH�Q���T�<Ar"Oxp�D�ވH�v�EI//�*L�p"O��c��C`�"���:�0ى"O`�s�߮'�2��Ǉ]�>ܐ�"O�����$d� ��P��sp
�*�"O
�)�m\�|?��J���]Y:U�"OJܲ�_Six+� ߔ=�h(YU"O�a)5n��"q�p7���"O�в�	!����A��)S"���"O0��C� a�0�H�H9">���"O]z�k��E֔DC#W$h�"O>���[+X.��0�"m��!4"O�r���3�P���b�����u"O��A��
�@�ȉ�WoѬ]��Ѣ3"O(���-ަ2ä��􋞀>~t�T"O�bH�,C����-µS��=ac"Oa�%��|����c�>�XxD"O8�;��T�b��{'Zy�D"OJ<�S�g��e�,Τl$��p"OR����<��yR��FV�d�"Oѳ7&T�_qJ1q���	D��੓"O\�K���#`��5)  �7�`���"O��rO����5�������aa"O>!��2K����F�&	��Da3"O��5dڣ(�4��d�)y%��"Oc�ݯVH�	Ja��.�X��"O~��'g\ ��Y�!��%f�0���"O~0�V�Yo�4�#N��~� "O�lr���a��Y� �>$�K�"O\ 2o
�z��ɰ���r�uy�"Oh)��:D�<��턋s��"O�9X��M./+��� ��v��!"O�q:�e��]p��p�A  ����"O"��׭p�Re�J0:�PP�"O�ĉ &��β��d�D�$�� "O��RV�^�q���"����*�"O�a���#�����I{>`y�"O�+I�Eղ�s�� 0�@"O��8��E [H�@�'��A|̀3"O��p��$����ꄨ� z�"O��z�肊 -<�	H#�&��"O&��ҠP�b�6�@�V�wC:|2"O2y���vG�qBN?$���"O�t�r�X�g�D���!ăsD {U*O@���$� U���ѠE��"�`�'�=9�L�Dn��v�{����
�'��1�.ڱ f�a8�$Ut/���
�'^ta����=�LtS@+=I��	�'O$�2FB�6b!L2Ee�9\�S�'�Y���u!N���L=F�L5
	�'�� �R		�
>TS3�ׅF�܈��'��觥��+�:�%Q�I��8��'��}�Q�N�K,�a�B"�Aǀ���'/����&;T���c�8"�
 ��'�>AH�OӌA�����c�%���� �ъ !+{g0Ԓ���J5�Q�6"O�����?��#'Þ*Z!,���"O����)�R}5��� ��Z "O��Ign5!6L��������"Oza��n6����o_#9�:\��"O��*�ͼq�$�����48��T��"Ob�Z�Ŋ^��3��Y/>|�"O�X�o��|��k�n1�-jV"O�ԱA�)u:���X�r0`@"Oi���$"C����ზ5U�!A"O�����R�K͠	��ec�%�y�&I�d|��� �� |5F����y2��v���`2ϵr�f��S�ߠ�yrM�rt�H#��+m.֘H�$��y������� bN��;�y"�p�4Q�F���^�d��W�ڽ�y�l�s[�}����A�8#"�ʻ�y"��wˌA���f��LH�+�yZ�p�p�`�c����l��Ȅȓ7�6b%�X�7�D��)N {����ȓ�@�Zf#�.h+������a��OǼ-Ҷ�R�jj��B��� b6�$�����B�� n������Y]d$���8�Y��"N 0�X��˭b?\���Q!���+��V.�m(��C�}�6A��>��Bp.؂8Di�d�
x`VM�ȓj�f�p�տ5w�ap���`��ن�sD�`��!e
����2wE��������N�!X�H�/<����i?�����F�R�[�L߅&��L��I��]"Ҡ]�?�8���T�
�ȓw���j�D�=C��q $�9T^��0�.]��G������GbY4'o`��=�ա k��IJ�H@�ï1����ȓ1dT)�AB�y����@�*7K�Ȇȓ{�z #I{�B�H�&Gp�ȓZ62
c��;&Y@Hv�	� хȓ��E���V�w�.iq�N_�]���a�5J�\>�	A�NY�l���ȓU��d��䔊p����˃ T`Єȓk�<%��#84HR����lń�K�n!���.M�D�5�Do��=�ȓ%������WԖ��Vi���Y�ȓH?�i
�+@��>����{2䱆�y���D�$\���MӲ`*:x��}_0q[3eG�)��$���I����ȓ((���BY!?"�*BFW'`�n�ȓ
�X!�#"�.Z_�E"��"Y3쐇ȓ^�J�1F,�y ���4n 
^�H�ȓ0^r{�j�D�Cπ�P�|��ȓ{Y@�m�"hj8=�.�3x��X��:�m`����I�6+ܹD����@�P7�؋)���Rh����u�ȓ؈+����Lb��(G��#~j��V�&�\�[�h[�c�9�����.a�]xdز79��X�x����ȓs8〈�E�=)7�)��`�*9:���JL����*0P���B�A��̅ȓ<�,�Qp�	��q�4%��~�Ĉ��SNL%���#��t�Sb˔'��=��ożqi�-��� ���"2���ȓG����U'X�X ,)�hM#��U��:��]H�HR�(i~�s�A�y}���R�,URwƁl���H1e��[�*���S�? ���,�!�v�9��� v�8�KR�<��	��FE���6�d9Xrf��
�B䉉L��Y��-O3_	%)f��YY�C��$$�L�e���Eĭ���=k~��D6ғ.��1��JB�E�F�J'Z�o�����i�y��#b�2qo�l����
G#D�d"�*	��	�Ʒz�!D�6D��Y�h��^5
��E"%
���8D�|��;�l��#��8Ws��蠪7D��* �X�
�MÑ�M�b�*7%6D�xb�*ܑk�d|�U��9eV�]���>D�F�@���/�0S՞E�Qc)D�,���[ ����Y	�H�2D�p���n;8�k�OL:B�X�*�0D��B��H�kԃՏ|�� ,D�lZ4���I�E�BT.y�B=���)D�h�@�& /�q�RlܜDAn0r!C'D���C�(?��`[��Y/_��K�n#D��y�/э{RxFK\���i<D�PB�j�8&��<�w.�8r��d[t$<D�[�N^*#B�H����9D�<��&[��Y"�,Y�E{~hӅ�6D��t�	3w��Q�$[_Ub����6D�)!A��|���`�
��JF�5D�(	�C�|�ӔJ�,�4 ��9D�����8_H<���O���i�F%D�pQ�̲s�QxD :KQ�S@�=D�3�)��I��u�"��a:��r�:D�q�A�:d��0�]+EO��Xf:��ȟ�p��ak,����X V��ۥ"O�@�q��laE���bf2آt"O���"�"=��lbWm��G+��f"O^���KA�?~�IK��/ $�+�"Oq�\"eYdD�WJ�m�ҥC�"O���[Ur}��; ��@��"O0��(jv�ŋQ��*K�X��"OPu{��ػH���l��xBA��"O���LK��8'�N ���"O´��J�/�p��c�;���zT"OP �įϞJ"�e��]�r�Ĺ�"On��b=2��͘���L�z�hD�>�	�7� 0�7hR�GEиc0@Qv�@��6����e��z�ĥ�v�Z2����ȓS�4��Wlߚz��鑨�D���ȓ�ĉ���G�T��	���dX(��ȓHDܠj@�ZN���U��AW�	��hO?�5��"��ЖmC--��V,%D�zv��8+�xC��,K�h8�u	#D�,�@#�OD��ɂ�!�,LJ� D����bH')���BRO];n��sv�=D��R��@�j:h P�1T�4q�<D��z��7Z{v�׵�(��">D����R)����!�S�=�EN1?�����7@����g�#a��D�*B+$�B�Ɍ)������ [<쵮�Z�"OƽH��
  ��A/�? ��g*O����B�vp�ǝw��}�/O��3�az�ԸyV<��l-� 8�Ϝ�yb�A�&�l[6�O�d�� *G��!�y2FM/-�F��A��
����A��y"�׌G��}@	�8|c�i�RGݔ�y2%ETʜM�PK
c�t�J��^$�ybI��/��`�]$$-�BfS��yb�7	�����&��\�F��!�ҝ�y
� �HD'T9S��ĳ
�b��90�"OJ1�f-�-$�����7l#a��"OR|��Θ9Y+���#(7�Lې"O6D�Сj��k0��B��!Cr�<I�i�|ܞI��mƀi�&�cP�\g�<Y`S�C���
A(� J'BM�͓{�<�Eǝ.�ڕ�O�e���
��]�<a�D]1y�npWgV�0��q6ˑ@�<YR,ָ	<����k��1�q��@�<Ɂ�_�i��TZsb�tz�<K��Ɵ�҆�')��K��ЀB��8Jr�Z�Rۦ�[�)�>�'׶�K��D�.�di�1炑w��1�'L�p�nօ�g�Ɍ�$9�S�4��>2��1�ƥVK�lBFω��yҏ�;m�����l�"G"|P��ē��y"��);|0� K�5P��Ip�K��y��� �Ѝw��>Lr�` 0�<�yb+/���B�7����G\#�y���/wmD�W1஘��O��yB�/j�VP�����L �@'�y���0Z����HH��n�Q�Z�yb�1��	A/R�~̰���y�aW:v�����l�JiP3ŏV��y�dB���T@�+K�D/|��w㌘�y�͏$Q�ܝc@�3O�Lу�O��yb@ڹs��	�7�&Si�q�%�;�yZY�h$�����-�E�V��fB䉚,LV���&b��:g$�{\6B�I9`�v��Ǆ:Y�Bɻ �ԓrB��69y{�E�L��P�:O8B�I�u>2��3�˾\�p�)K�`$B�	� h�;A���\��|�k�>K�
B�ɽ~���C+�s���Z�	��C䉯$��Dx#jO2ib��3����`B�I$0��]"�<L���hGd^%ENB����RK�h�\șܬ�<B�I�UD���G�O�$Jhݢ$��5"O^�0F�OCq��q�̝/��!�"O��0�b�'�E�cd]
AQt�8�"O H�cf*k2ȸxB����I�"O
���5}$дH�n��e"O�t/BG�ɣPN�>e�$�"OX��UCDO*]ꦂ������"O\I���!�a�H�CބX�0"Oti�Н����`��u�,9�"O��BeA&L*A�{j����"O����O:8����&��(E^$Qy�"O��Ӥ�+�t���+�ZJ�H�"O6�pq�٩"�"��ɔ�JTLI�"O>��k��$E�0�H�m��m#t"OB !���U:�(9�Y�^���#"O����&^*)���.|�(�k�"O�	���N|Pp;6$S�r� h��"O�I)�eI�jmDT�eջ�d�@6"O8$���P(+�Z����E�\N�8�"O0��D�5V+�(�e`� I��{�"Ob��C���7s�K��J�S�P��"O���@�Ъc5���nG�F�4M��"O�DbFŉF	�t�����M	�"O��9b���!��(rJѥ�j}h�"O�I�R-�4:IѢ�0?p�V"O�y�(|��d���قnk�X
�"O��;*�3f�(�2 @	~ ���"O0���&R�0�����,��0v�tQa"O� pɧ���mch���Kˇor�т�"O tA�M�2k"�#È	�%j�d�"O�d�q��+,�Pp8�gsF��p"O2���e��J�ƍp3@�*56���"O:I�0aR�w���E�٬����"O���B����p#t�f"O����,\�,�q�#�5vs�E�"O8m�#Ѕ)�h큲%� ]Z�T�p"O�A �Ƒߐ��&% �rW4]b1"O.,�֊R���*��P�F$Ʊh�"O��Q�4C=rx��b	�rb��"Ox��@D�%$k,$8⎿~��c�"Oܼ�U�	EIP��'�	�ex�"O&�����xl��ܒW F	!�"O��2�A7ܒ= ������"O�l���H�e8١5��H��"O�L��gP6>�\�����T�R��b"O qhw
)R(�4ɜ��t<�"O�$�!�"_�!3��Q�m˪�:�"O������hM`a+!
�[h�Dac"O.H`�!V38QN�
�ɓ�~^&�B"ODbV��~�2��#D@f(�"O����E�v�ؼ�b&���	"O��s㔹DόY{��Ȓ<�T��v"O���[�Z�h����1�0�B�"OB=Y���T�����H�e�D"O�4���)F�x%��^�|�"O�<�jTXl4"��!S*���"O�<8W'ݘ+Ӝ{d���u7���g"OTP1��#p�})&�Kd@b��c"O�e�X9�R��@)�B�p6"O�"o��c�HL1Ce��D�ĭ��"O�ᆫ�jf� "���'`�& r�"O�a&�T;����!B=x��8(B"O�-seAþ!�\eÎ�`��1�1"O��)V"��p>��я�[����"O��K`/�<��9X' &:��"O��HJ�3\�W�/We�uۅ"O(ZVv���B4 P�vv� 3"O���D*��c�[���R�"O�M
�j�<Y�|��B�	� ��"O�xQ���İ��GK�d���"Ojm���	�\l�Se{�&�0@"O�ɀ]p�-��Ϋ"ńA�"O~L�f٥�b4�U�Ϩ9��q"O�]0��V,��`�B<}�ܘf"Ox���M�v�@	� �;"$��"O�R�-X5$0�t�q1��"O�Q�$'H�{���r�.N6�$�3T"O��s���O&�m�	���+�"O�����Ũ$���e��� t��A0"O�5bC�&,�=�d
W- `��K0"O~�z�
.`{4qr0�#P�5�d"O,��W�|0����eo�!1P"O^8�RAG)� �2C��'JDpE;�"O4p����D6���O��R�0�"O2�Z�������2���-�JU�V"O��(�]�B}q6`MY�`�$"O>ոčK2`�7@�,(���p�"O�A�bAV�q�MA�'yq��q�"O���ҋM�;��q(���j����"O�Mc�X�i�p����p�����"O\d�'�5��lI@H�.����b"O�IK�/C��}���P���"O� 4�  FN:n�\��p�O>c��"O-�%^!� MJJlz����"O��W�B%�T v
J�`x�(;�"O�-�vc��֜y	��(d�R�"OZ �c�5B��� ��B�i��"OޘP%�$z���C(�M��1�0"O� r���:?�Ƚ��&�&�h�#f"O�����>~�x����m�����"O~��0`�Fb֨��	�w����W"O����M@�rh����.)h��&"O��!3�� B�X�]Iܴ��"O<����
�j���g�ꭳ"O��3RC۴m��K�NC;=]\�`�"O���D���< f �TNV<oW���W"OYz�e�4d��B �Ju5"O`�ؐ+�-�j�)�o��zF8�Xp"Ofz�i�0{��`8wE��chY�"O.�Rs��)n�2���$��ii�"O$�3�F8�R�)���q�!*"O�Yqm� x�����'�^8�%"O�Ub���;X��HRե]j��h�6"O�]cg"DR�e�eeO�-ބ��"O���U��um�p��4%���E"Oƌ��_��Ts�E�2��t0�"O�=i��߈P�r}����~�|���"O@L�4�ض���9�n[���"O2a����>o���rn^]xx�B"O&XA"��n;�)
b��
ou�РQ"ObY��-x�P�1怓24gx�Q�"O�M�b+�M0�MC�otp�a��"O�@��˘lh�U��nz�Å�bq!�DN�|x๓�����x�d�&Gk!򤂅O^���J�X�D̐)�eS!�d�5}�����̽=����&h]?3@!�D&����M\�����؎+*!��B�ჰ�<s��lS��S%.C!�$��R�u�&
2�Đ#��БF$!򄄱7`6P�"X�٠��B�n3!�dQ��T�"��	r�Ha H]59!�ZOz���띂����  l{!�D��#\(+�k-�!�7�ڤB�!�H�k��(��E�����3�!�d��	ᔹط.X4s���U�-[�!��G�&\(�a�7i��H��ڀK�!�1K?�9b����l��� �!�D�hm#U� �=��a�gEG!���4w^ܫp��T�B(bRl��x!�9�k�,H<Q2@��RQ�!��Q�Nv�Hw,��X�`� Ti!�ջ_�8h�g��f#���a�+S!�$S�%YZi�s���t���D!�$G(p|rV�\^ L��q��*~!���.%��e`�EB��C�L��mi!�A�e���[��T�EX@H��ܟT!�d
�zk�����"�j��4�S�~V!�d�� B6�	a���}��D�!M��\�!��]�&�ڭ��A�+o��pU�Y
!��%��I%%�NG�1fµq�!��N�G���a�)RC��t��7J�!�
�Q#NƬʜw�p����>�!�����pЄ��\ �P����U�!���.|�,�7.R �,eqD*$)�!�V`�qh�Ƒ9�N��Ԉ��v!��L��&��! ���<PЦ`!�� 
9�h�-`dD� �O�dU
��6"O*�A�i��fc�8��%#tQD#"OJ��wJ\,t5��b#{=�l��"O�A��4\㴅iU!O?&�,�"O��@P�(�\�X�O��7+F�{�"Of�r��??�^;3�E�s|�Y&"O�C�iǊo�^�:A����:V"O\H��
�;TL�XvĂ�s�ơ��"O��!d�<7��l{�m�;��xF"ODD�e�>\1A�K
^QB}	�"O� +��}늩�!k�MN�S�"O(E��,)M7��o�rHn|bv"OT�@�m�Lx٢q� �y�"On�v+ɲE��)��W!tF�)�V"O`u�`�W�D�0�0�5QY�D!V"Ox9:��1Y��x�!�C�C���"O8�P�hR�+@�`q�d"O�=��cZ�s~4��D<d�$�"OV�v�ǵjJ$mYW����p�"O���H,�>a�ԡ�8}\#�"Ob�;���Z���/U�%�P��y"�K� ��r͏�ټ�@҅���y���������W�a9�	�(�y�n�>�f�A$��0�R
RGP��y"�O�X8�[��2~3�@��yR�Ƒt������vº�cC�V�y��I�diև�!g����G�ׅ�y�*��C�J�k &Y	Ju'%�,�y��
�2� '+�P�ܭ��DF��y�gĎ���p	��0Ģ���E��y�d�<-i��;���/�N1�w�J�yRb�I����2,��[#��&�ƥ�y��J%e��h����)-e�����y℈5uR4�ࢤ�i@.��5���y��M�n+�lq���b��T��U��yr�e?� kfhǏg� �C4!
$�yrF=}�(�`����o�FM������y�B�3~�tX��m��؄��yb��N��8��F�\�4�+��%�y2��"p�@EY#\qZ�6���y�)��"p��чC�0V3�qJ�/^��y���5 �j��TÞ�D����e�_��y��#8X�B�-��B2���ք�y�)о?m��Q�M�J��`dFK8�y"C�|�A��'sv\�m�y���m'(�1��o���"Ä��y U�kb@�i��ݡ3[r�r�ç�yBo�Za��R���v4|x�Tf��yR%E?T8�lٗ"0v�����D��y�������(M�u�Z�A4�M��yBąT �P�gFO�A`$������y�G�*�ܬH0D^-cW�&B��B�ɛ�YK��H�X"���pI�:$fB�ɢMn� �ĩ�!15�M)d̚RB�ɷs{N���Hz�y��ڦ�C��gx�@Q�܂!�@%�7/ֈ�B�I9G��t�c
G�.��4&R��B�I/βؑU�>*�ذ���3a`B�HHt�Sf	/[���-N<Yi:B�	?EF�E�ǩJW�ԑѥǽ.� B�	�kt>�+'h���t��J�%J�HB�I�+�
Qa���)�V���j��e�B��+�>8RQ�
ALLR��(�C��2!J	�v�[(-.0��G]�
�C�)� �}AA�)3\,E8��5���"O^�3��I	���;G&�.-�,��"O�I: ���`�]���L�/%�p�64���f=Nh�\��#� �* !9D�p�p��n���Ae�)F X���;D�`qR����LCr�M	,$؅�?D��k�`�j|��V �dz�A=D�d9�&(ˌL����X�~����<D�����.�0-c�Q�t�PXՌ<D�����/�𕊳-�_`QC�$D���Pύ�"wp��8���!D�d G]�v<^9�en
�2�88B��*D��ѷ�Q�ELԨ �,]�]� �g�3D��p��Q�+�䄁�AE9����J0D�X����'ZX����Ձ$�8D�tS��!�nT�ϦeS��q�$D�Dӕ��/�,���o%���2n!D���
Lˈ4�5O�&(��9��:D�L*sDA�q�~8��`.��S��<D��8c�PO���L�/R�d
9D�����[ ��U��9ڀ�	��$D�\��G�Z�>9�-A|���B�7D�؃��{�Bj&)�1C*��pU�6����OW��Q ��
� 0+ဆ<_v����O|Ś�Ǧj�q�3a�,W�tAd"O��I#n$'_����	z�t�a<D��SE$Y�(\����|7���i.D�$����h7ޤ!�*�R԰´�/D�x�׮��t���ƏD�
����(D�lkG"��?��B���' Z�#@1D�Pࠣπ`~�Qؒ��H�t`�+0D�`����(: +��+
�
x��A/D�t�!��$�X�n��:�,�&�-D�T�����xU��M`9I%�.D�hrӂ�6?���:��Ix��T�aM,D���p-W�5`h@�a-+��$!Ch>D�TCH�N���+��S  �����(D�|@�	�`�PkcC�=l��8#��(D�̚�NC�Tɞ4c"A�W��d���2D��:2K?�ɻ�U_p��a,D�L���ҫ��#vF�!S;J1��>D���v��-zH����!�(}��0D�
�#j��P�1��
e�X�S�(D��K$�9:,�c��*��נ(���&%9��������AP�h�)I�"Oi(%DQ	Gj�* ��\`\��"O�U+!#�����e'5�d�z�"OBM��C�I�������4�ܰ�"O�9#��M�%��1"�" �  �"O:��sDD�,���iP�x�"O�u���56��x�G����H27"Ol|��l�7	�8r����2�&ĸ�"O��ó�Y�r�,��X3d�ې"O慁v�G�K� a��խ&�k�"O�Dyf�'^e�2&C&e8��"O ��b�֊������;{��ْ"O6��!!�<tw�!�B>{H��R�"O��g�|@D���DS�hY�咅O��$��D���I�77��;���}�C�ɶK	�� �n!�h���I�[�|B�	�J\X�dǢ%���[�izr*1D�P�uF.�F�׌H�=�p{�3D�����F&Ee���C�F*a����"l3D���V�:8���s�
!j�4L0D�� �s��0uX�MCDI��^ٙ��'��OF��a��m��3�`E�Z�$;c"OV�+�]�LJRM�ҏ$���Zp"O�HX�X�LH
�H����8z�"O�mF1�$��B�ox�yZ2"O�4�2bK^<�)D �dՄ0��"O���ԯ|�t0�M����<ҳ"O��qvI^K1c�F�Z��X��'4�'��]� ��4TFL$C�`�l%1�'��0V�L�Rp�&�QA\ɒ�';6�#�l�/-(���ƤQx�1
�'KJ���D�%�2x�׾`E�P��'�Q�ǞL��Pi�*�T'�̠�'xm����8�|�c�� ���'���4G.Ez�����vf��)�'w`�3�:�d]�R�еsӴYj�'��s�⇼��9ね�m��`9�'|,P��*gÎ�a%i��;�'���iZ�v�E�G�Ʈ^�M��';z�31�����걌K�P�4�y�'d��д%�E��ԑ ��I�' 
�@!/d��m��!ɐg�R-�
�'@�x���� ���ת���vк	�'y0��O�#l� �V'ڕ<�H��'|`YR�Ő��l��%�>.m0 *�'.�T�e+�8��{��6%�`��'��	�@�q�\@{$���$��
�'��H�a�6AxY`aĀ�p�U�	�'#���d�4�zʠ��:o����y��)�S���] �jH�u~^�0B�ɱ& �%��!(�6d`G�!=�C�ɉ}��@���ie�K�@ML��C�	��<��G�Ѕ����l�B䉦=����Qk֩C���;������B�	�X�ֹ�$Z�C���b'J$ A�B��U������H���#�Rpz�B��.<��&MV���r�f�Z��C䉻JF��pcf<X���j��I]|C��
4��(`j��	o���QH]gRC�I�MX~ĺ���yv�S��z@C䉚YYؼ�p�	?���0@,�#+C�I�o!$9�-���yŋ��B�	����Fɔ'Ċ�CEό���C�I�7�va�$�ҿfJp)��_ >��C�	�o9�ݹ�c�͆�
q�E$b�0��ȓR�j���N�0BG$R �B"W����o��L
c晠F�v�4���|䜄�E�
���Ҏ
D����EE�0��ȓJS��!2�O����.�!jںL���� �C$I| �t�˟1��h�'��}�j����hK�K�$W�X1��P��y���qh�٧��L	*e)�gU��y���
N�( ��
�/J�ܑA��yB��|�E�]+B��(��[��y"EѲ�PKb�<���ϑ�yN\�g�4b�"�:x�������0>�I>Y�G��3��,BG9��dزG�<	��O�yҤ��#]���2�^D�<����{��5p��>��;R��<���bh�X� ��n�җ��}�<	��]�.�P���
w�~�� q�<9¥��k��8��Nl��!�T l�<9S.N��X:�KG��n���Ia��@�'����'(Q^�؉� N'ҽ�
��� ±���	7� 0�`��rA:q9�"OЉ1$牸j�vSemF�0j�1"O��{囜f��;`
&�$�"O|%
"��4*���M-~,]��"OԐ8�n��yغ�˖G�3d��M�"O����$N��%��͕~��t8��'��O�E�tL�<t�س��,M�np0FL<�S��y��ЬE�l��r/0'�3�0�y8{hz���:@X�v�ҧ�yB��>!�����OɑM�����T4�y��[�lb���+\��96�ɚ�y���r{��Kqj:V����Ĕ��y��P�#=2TA��J8��:�#<�,O:�}��nȍ4�\�"�bq���R/@w~��Im�	�FL"��b$�!��P�Kܜiq�B��6G�4��!��>-V�4�Y#��B�4L�X�EEw��-"1횋oMfB�I4�:A
�
V�#$b[�jMbB�	j� E�Gh��g�����$IxB�I�{W��Q����?���+� 
O�JB�I,ݖ@S3��tS�L:�f�>�(B��**:U`ƣ�Z^���"ً��B��,H�du��#F�~�8��	��B�)Z���'�ΏUz�4�'��>�B�I�G���u&D=�B(E/ϋk�zB�I�\�lấ%@31����0F�?!B�ɼJ�Z%� �3��0{7(|��C�ɠX+"MʀȊ2�����@�*R�C��jB���THA9kþ�{wꞋ�JC�I�E21�P*�X��qgɣDC�	$�e�Ə�JF`D�J�p޺C�ɖF(F���� Z u��Glz�C�	�D
�[�-,*K���G�o.�B��""�P��C�3��UYF�T���B�	p[����4����ԄK��b�,E{��D���؆� f^�F�9
� E��y��o��{a��M����/�y��VT&�[��y�R�����y�J��yy�ݺ*X�@3�ɱC(���y��ͧ'��pRe�m��P�C�"�yB��-[`�9�ĎmR�q	��U��yb.�G'H	�%�7V�qp),�y�#��DZ����u�P&��
�j�ȓ �i(E�7��mq�a�.�(q�ȓdn(3�A�5I��AՔZ�E��4�z�s7螏6����;G���M.�&N8b)���`��^��	�*�Sq�C���P%�Ň�jL��&%�·62�l̋�����ȓY~��s�Q[��ȣթ�aX	��#iȱ�v�'\Njy�'M�C���ȓQhA�L܁��RbU&=l�|�ȓQ# k!�8�@)�q,��{�v��G���1.�V5��QjPpTH��/�Z�AF�V�1�v�Ȣ
�DfN}��].�T
C��3�Ը���2(��?����B�tW�ܰ��4a{^� ׏�b(!��;A��`omhUCWl�=(!򄂄���!��"~���y�͆�!� 2x?���bҮZU�  ��L�!��.[��8KՇԕe���z���H!��7�l�p)�{9��Rf��&�!�ޗB���j�r����F�$S!�$�gt�3( �M��q�2��U0!�� .�AR⏷HJ�I*����	�"O�݀�ϡp=ʌ�k��3��"O����w8yȶ*\�V�c�"O�� A;����i21!��"O�y���G�m�r[���n$>}K�'��Ou�a�U�!�r�9ł{�Ј�5�ŞIi���x%��0���ZV���ȓJ�,:���+N��0B'ީYr����r�
	�w��	k�^�C5��&3ȍ���01[  �! U#��V	�\d���d�dY/iWZ݂���kfB�	�h2MC�gE)C@��d�
(s�">����ȋ> |�cᄶs���3�B��q�!�$�n*�t��j^�E�Bp2��s9!��'i��(��%��TӘA
�̕s!��
C��XI�mד�����	�.�!��]�xq�@O�
��AK�K��z�!�dţ �;4Ɋ~��iᵄ֌�!�d��/�����T��!��#��!�D��;�|�P�PB"Bq����|"1O���
>'0�3����L~V=Bp�Ĭ3;!�d�Y�p�1�@$gv�<{Tf?!�Dy���spF���p��:e!�d�R���Ф/�'���S7@Y�!�d�-����!�,{lݢ�(kb!��^�w4�*rM��D\z]�a 1Z!�Ă081�m�R���qVda�w�
=N�H��I�se~a���a%B�!�h̊z9zB�	ne� �l\�;'V,s���|bB�ɢ.�\r��B ��[��^�9�`B�I0?�������
����A�B�B��Z�Q{�$�r�.���͞�8<,B��t���(��$a�H�� G@� B�	�j"�9ptǍ�v4���%?B��mv^�Z�cW4?��ՁX�!��C�	�*�3�Η����˔	_�C�	�����u�D0*z� �*��(�C� �B�kT�	�m��|	��¼1��C�Iw��D� �P,(���`��C䉧w�T�8����V���)�ZC�I�Q:�S�,^�w�aB� �NC䉂l�H}	�n����`g�~�(C�ɔyJYQe"��02��A�I>�6B�	�
17&�"�s$,Z��DC�	�bP�j`���+��ԱiD�DnC�	`���E
�}�|���� �C��lAfs�FȺl�p�Q���R��"<a��4���$��m�I �_� 2��c�3)�1OH�=�|��R,oZU`Aė�I�օ���Yo�<���CI{J��1Eϭbm̡���g�<1��1[��;�M���D��W�<���!��Hz���$$�S�LR�<	3�_�����E�'q���J�C�<q��mx���`�9�A����B�<qbQ�V-�J�3VS��#�H�I̓��=�ǃ=�4ؗ�7�4`Q�z�<�0X>i�D��J71u|PB�!�K�<���.H��j2��58�(tz�c�F�<��Y,~4\rR`J4GÐ,����@�<yP��?AZ�
#l�.Rʠ8����~�<ѳ�ϙ/Z2����h�T�����`��<��؟ p%�#H�A/ǁ3d�1(�:D��1��7,�h�X��ŉ��]sd�%D��֍N(c��uK���H�yQ�!'D�� @�B坚�(����7	��Ő�"O�����״���pu`��F@2��"O8x��l��x�t��D`ލm/:��#"OBh����+����H5]���"O�90�!|pԹ	�n�	�2�a�"O`�Y�k
֤�q�g�/|�^�Q"Op�qtF� �Hm����`Cf	�C"Oa���ܷNXI�����J(*�bE"O���	��|
��u`O.<�H�"O�|�r��-_\<�����/�<0`b"O����P6(?b�:V�I��
�H2"O�̩bI�ᖐRQ*ڰo�Dx�p"O,Yz#�0#��)�gџ>rjA!�"O�Xr�j�?dč�w�
�3�P��P"O,�R�A�>�D��A�D� ��"O>�xSNѢ|��Q�없]Б"O��1&��m����*[�Wg0%Ke"O� ��¹qS�������Il��"O�@b���6=�
�
F*�57b0]�#�������dg�`E��,��qB'G	�}7:C�I'|���3�¿ ,�)��3 
C䉗^�ÅףB;ņyk֤��T2B��?"�L����*$�PaRG�B�B�	3\�̩�c�EY:�E���B�	%}�$d�} Ab!f��,b�B�I�r��y��� b��DV�~����]y��'�>M����[������T��u �'l��b��W;(����'�0A4-X�'~pBR�#\l�hp��޻<��X�	�'G�@Sǎ/*�x	v�N55x���'��%��3a�a��k�#�H=��'�,���Nr���2��O�����'})���\Izt��� ���'�R�'��{B�-H��i��,4EQ����Ѐ�y�e@+��yb��B\�Lڀ��y�!G���l����K?Z) $�(��'z�{b�1[�k���$8'F�#���yԦ"`���bFN�7(Ij&�:�y��3I�t}+���Xs���I�1�y��S�"8������z���ө��y�"W2Ӱ)i�i�H)�Pb�H͝�y"�ߎ? �ZVRl��J�����y�B9Sײ�*e�u�"�� "͍���;�O:EY5I�5T��9�o΃e�z��q"O�Q�坙NR ׬_�n�ڝ�"O8`��F�QT�1���T�6@�e"O$t��(M"y��@��A
)��uyp"O�%����QnZ�3�G\����W"O���kS��QZ��'r��(��"O|�UEݬ@����D�
���#�"O@�0�	
	0PQӗE�M�ޝ8�"OH�9#N>$�֔�e�p�BI2T"O��#�H#:�Z���n�(PǴ9y"O��e�W>vH���dxy�"O�ȑC�*4��X�D�ݍzM��ya"O�l��C�,�<�³(ѱ{YLS6"O!ʇnY8�t�i��D W�
�"OT�����? ����\�W
�x "O`�ˡ�˛<��U��գHV0�B%"O|y�'G<K��U����.PVʝ8�"OF�tK67�9z�@L*7E�5pa"O�xZ��9�Ң��N �*R"O.��Y-4,(qA=_	�M�"OZpC�I�K�}
�*����"O� :Q��Ȟ%?$�%ڠ#J�*8�"O\�J�m�lʖ� �'�O\�W"O4$��cC�R�,�����\�*ش"O�E3D�Ԯ{xT��g��*q�6 ��"OV C1��$�pM��^1IHLU�`"O�0���ʴN
<ix�B``"O.xI`�E9x)�)3v�z��`)V"ON��ABA:O���r���@L��"O�$蒁̣Et���̀ISlA"Ox`$�H�K`���(��$���e"OF9j#��<(�1���C4�Z�"O��hDǙl&�a�fF�`�5��"O�H�4��;��}+C�Z��3D�H�Q{b$�ȱw-�����0D� Rצ�o��p��%e��`�2D�����߭2���A��wC�P��3D�ᰍ�)�>�Y��J<�|��%E1D��H��/jQ8L�F�K�Y�L��Ј!D�䅙w�l �'i��f�p�r�) D�K��ޓj�,���B'R�R�>D�H@@��fƘq7B
�"���1?Y����i�	EÃ�+lnQae��nC䉦t�E�PIH��`QGg'\��B�	����:��I(����0��x*z��� ���+��ER�h֘Y��p ��z��	{y�'�8,�7 T<e�©(S�N匱��'h�y(�ұ;�"a���д
9��`�'d��QG!�"@��è��:
�'Mb���o��/�����e"]�
�'�Ĳc�^+f��0e�b��'s�X�I��jp(- �k�)O��h[
�'�F�ɀA���0P�X5Rs�9��y"�':"�Z��1=�(|�'"�&GI��B�'I��9���Q>��榁�D�Ƚ�
�'��8�����%g�@Sn�8C^Jp[��)��<Y�/B��D �!��j�Bx��!G�<��W�=�P"��D�P�c$h�E�<��/\>�ڰ����bzh$���B�<��hyI����H2,�$J(0��#>�-O4�?�많�=tE �á�F����� D����`�	j��r���%>I���:D�䫑EZcl�q�0&��6���Wr�����$ι=�P��c�Җ9UlīgO��!��S!J.�}��"'?H(}ӎĐj!�D�=$�d���9�ԛB��!��Tw�]�"��"�U��䂝k�!�#:zt���e�S�\;_�!�D[+I�n�1�H��N\��b��	Yvaz��T�/p<��s(�!L�܉j� �3r��'�'?=��(Rx 6	�b�H�9�,D� �Fdو_�ZȠ�V�/0��D�*D� � bژml%S�KB]<�ɧ�3D�cpץ/) ����0廣e?D����X�(���Ɇ�^�{��Ja�;��hO�S��:Q���v��	�5'�5H�pB�I�LdZA@T�L
1�A$%�Db��E{��T�e$�I��G[2 ٸB���y⮐�)�@]�oN! ���Z��.�y�%Zd��kC��>b��J�x��'�u{i�*�@(
ԏ�3����'8��TfE�S��x&�I�"e���Ox�=E�d�U�Blt K\\�ҬQ���y��)�����9h�"Q�1%	�7T��u��z�<ᒊ�9�h�dկ^Enm@���<� p�bv�ɥG���6�ߪ��hC�"Ob��A�YMBY���t�Đ@w"O�ـ���-3���QCO[��m[2"O��!�j�"P���pO)� AS2�	|������u��'�n��0`��"#!���OX�� �B}Q���h��r"OB��'�V#Q�5�V�=8�p��9|O�U�v��(�N%����@�j�kQ"O҉�.\g����&%�H��"O>�pE�^�)	��t�-`�yyq"O�c��&T!xB�	�l A2O���d�T��(��h�s�*!��j��D/�S�O{d�c��׫>) -)��٭LPE��''�A��)'��M����I�� ��'vt ��8h��1b�oX�p��'�ZL�'��(l��ma�b_Ķ@�'�H`p�Y�mں���D����*	�'ܮ4�Oĭ��	獏8ep�|���'��	ky|ʟ�d�� ,H(���;0�L���Z6'!�$�R�0��S�+0��%�u�!�$;u��jG�V���h�:4*!��U+D�D�8���
cq�5��h�!�$�I{>}�!�D@Ua���)!�D�*�4E�QhM��8ׁ�
%�!�Ջ;�>H��@��X,����^+F�C�9�Ī�.Ƴ'P8Ri��pV�o���2"jNJ��ء���P�T4��nyғ|B�'_��$t%V�
�2Bڄx1ۘIg!�_2R0���P#޺S���8 �?lN!�D�����I�<<�"N��,E!����qYS:���-EX7!�$M�k{�yG�0y*�����?q�a||��'J���&�u������y�g�&MQ����mh(�A��4��$5�S�O��T��~�0!6�-��x��'"�ۣ�E�56�����!�)��'�j���(M�+s�TK0��"k4���'��z#�ʱ?�ظB)�t�2�'��b�
?12$9d�1�,� �	!�0=�b�K3��Q��7��+ �,��'�ў�'���T�j� D)h� B��p�B#D��zb�0LL���F�b0�Ty�$D���䭏4R��+Ĩd�\@��#D�p��ĿA��Q�G-�7��P�qc"D�P���<�N�!�ɍ(�FP@�++D�T3r��;
�9��G�丐�$D�T���ց:���7��<�bd-��<��$O���
�͐/;��Dy5k[[�<���?��{���!_b���U/]}�<�qKS8u����@oZe�0�`E�<�'�X2Y;Pd���
�ꀺ!�@�<��J/i#��3H��m
Q+C�<y��0]j�`�.BLh���&�y�<����/�ZW�$�r�)�h�s~��'~L�i<D�&\ct7� q����<F�Ƙ;p�m�ۆ/2	�!�r�8�$@K�F�rp�P�7H�!��Pz형٦*:[��Q32`��!��ι[�r�J�K)�*���nE/�!���-I� � -��{������?�!�dƻ��i�`��h~0�@J�e�!��ɞT��Q$�6gO�%�G�4?*!������w�-=�`,3kE�!��P�U�L���޽a}@�SV�JC�)� ���ԉB;-�m�UG£���"Od]rWl���(U:e��eFPMc�"On	*�,2�y:O1>',Yx1"Oh�Z4#�B�@1pN�~P�`"Opc��K}x��S�C�&�I "O�x@G��Y�[A���O����"Oz8P���	ЖK5�C,�4`"O.٥��x�;4#U�lb X6"O޼��ɩ@� ��!	
<�BiX�"O����5�0ћ��+�0�a"Oa)�1M�^��� r��83T"O� ��#R�% (,!!ON����"O>=��cZZ�(��C��B�\�`C"Or�c�$'��`J�h�=� �	�"Oy�"�{�FU�g$)���'"O"᪡e���1�b�ǫ:ސ8� "O�q�#�=%�D8Ƅ*3ql�xC"O�Q�፳GdLl�-��MZМ�V"O�zF�)� �i��XDK*e��"O�dȥ*�u��#�,^#Rx���"O�D��.T�]�a0Ƭ�2:
0�P"O�L��o_(�4�ڠXQ>�V�>D�|��� ;�`\&/��'�jp[3�;D�`���\U%0�!���X�2��,:D�4c�O7pr����F[vT�2��9D�`���?T��[����
ALq��I8D����* ��k����F�Ƃ"D���)��d�lW��	�`�!D�H-\H�G�W�nU����2m?LC��fO����M�M�5# �
OpC�)]�B@�Dh�mv� �J�H`�B䉪"k��!�@Cܘ���k�#�B������+�r��K�턷S�<C���16���
�xK��0K�B�ɬLZ�m3����Z�p� mѻ%��C�I�d�0`	�H.T�!����6C���b����#j"�	b�C�	�,Mp�Cr�]�8�,���;;��B�I)g=<��拞C�
b��o��B�	2rb�ة�b�n�����T�J�nC�ɡUq�kG�ʂm�$"�C�.F�vB��9z�1���-_cL�(�AK	�TB�I�3����C'fV��"LB�I� ��$�ԫ}�, �"m�k.&B�=���0�P�n+hI$��Z: B�	+x�ݩ�
Бa���r��Y�@�B��q``y��*ݮL�P���o��J��C��01N��hR��B�����9`8C�I�(Ͱ�X�M>NMY�T��B�I�T	sQ��U\`��U*$rC�I)h��K�;>��ɪ!i�xB�	=>�X!�+\�1��3����I7�C��.K#�!A��Z?�樱v�C(��C�I3n\��B��T@Q����-��WlC�� 
]���AF�� i��0CdݒR0�C䉈'2vAs�'�gԁ��Y:z��C�ɢ_�u���|��j��փ;�B�	�|}��j%��0MJXCQo��dB�	>��4�0�>_��C�O�
Z?&B�	�N2f�a픍G<X��
X�B� D�,S�!M)21��#I�4aJ9c3M)D�@�䌕���)�ǻ5�Ԍ���'D���U��`��(��IW'��+��$D�Dȱ 
�rB\��	�q���3�>D�� )"��1f���'$�2!1��"O�ܘ��N�@^h[-X�V-��`W"Or�)������FK�a2A�"OZ5B��K��>I����2:���"O��`H�l��� ǖt�A)a"O>�
��ۦ.�D�'.I p��"O(Lrd�N�(}�CT1Q��9��"O����+9s��`�P	'���8"O �/A�1��}��RN��E"O���)�/97����cN4x��L22"O�� �: p�PK��)�Zd��"O����4���²c�����)�"O&�C`�4Fk�C3�K v��D[d"O&qH�bӖ+���,�a��`�g"O�t#�N'	
�ݒQM�0�`��f"O���� �Q�r`���G<Qk���`"O^ŰwA�, �Ce.�\���ba"O��h��S芵�퐏-�<�8�"O�䐇�w�H���K=%?���"O���/ D��*�
]�>d!"O�ȗ�ǃK/B�S���o̔�""Or1���Ԑl���1����R�$"O��ш��6�i3�'�ܚ"Ol�!�¨*�qs Gܻ9��8�"O���D�͇=m�@� -=�"O�� w��9/��P���@3F�3q"O��y�J�,K���zrL��L@T�s"Od��P��oH~]��w�0s"ON)�Q������1���1���u"OΥ��$�ܜ�6F�\B|�p"O:�y� ^#@A�煑%2̌Ȣ"Oz0�p���Y*�c��� N�ᓵ"O�:��� �;�C�1V��p�"O�T	�B�.�l��P�D�A���s"OJ�S�"����tZTċ!-
�+"O�}p&�V
$cEA�"t�!"O���AΉI�h��!K��N�x���"O�z���.&L1���O�!{��Y�"O�pbd"T%MR Pb�OYo0Y�"O����F�7*����o�+X��C"O�`ӡb���
e#'iP�S��D"Ol̓�m�<4��K�Aex��"O���PQ��^ـ�U�4_@&"Ot]����B���;c �-UBV��"OJMi�& 2lJ��R�=,4�4�a"OڤC4GU�/[|M[��³�x�"O�D�F 03�M���/�܀f"OL�p��w���Ä.��e"OR����ӨS�M��k٠c�~Y�S"O^�s�L
���`s��03��u�"Oڜ	A��3Vr<���Ý\�l���"O��� �9x�QK�j¦V%bd�"O�|���,wg����
MZ����b"O�$x�ʝ6dڍ¢���.�SR"O�:��X���D�Eˑ2��rq"O(�IP�69�.�!�Ő�B%���"O,�[�ήoe^�0��V$�!"O�Y�F8@�h�JC
J�H�F2"Ov��!C��{�k2$�+:9�!"O�H�D苻 qV�Da=���"O�@o6O�$i�&@@t���C%D�$��,M�:�R=�Ŧ��Z� 	� D�p{����~R8��![�P��H�=D��A��SU��+"Í�M8R�;D�� ���u�7t��}JS�Ů[��8��"Od"1`ٿ/�x�X�#�%RQ��&"O�`�6�v\n� #�t�xA�3"OZ�x�'�6�&U)���Kw��"OL�F�J1�A��܇vĺ�"OP���ǠT�:A;Gϓ#pjѸ�"Ohbb$�U��D�ˍ�nH���"OXՐ���Q7,����YR��"O걓�c@5��pi�!:;>EC�"O��V�R�L^A	�H�'o"��x$"O&X*��F���(W�po�� "O0��K�mh��[��	VS�%S�"O���/=|�,D����e�`��"O�ussN� CXN(V&�l�|ԡ�"O�Y��= N��c��P�"OB)0� �� ��E��ڙ 	��c"O`�����e�`��ơ����5�q"Oԉ�@�8��QbC;AS�m�"O �bJ=�,=��B��M��)b"O:R� \<|�@M�I�6aK#"On�R��3I���xc1q�
i٢"O�����w;���S�3B���j�"O��cd_[����!O�6�.� "O�MS6G�cP]���D�S�`8�7"O2��U���6���`T+W��ɁF"O �1H�m�ޠ�p-�-n��q"Ov���J��6���Dm�x���"O^ܢv�Q�nS��[�L�	.�Hݐ�"OE�E�Z�H�Pq�\2,�"�:""O�|�QeU���(v�3�n���"O����S<񒽱P��Y��Aق"O@!0E�J�����!z1��k�"O.�D	r�����̙*(��-a�"OE��H6h@{cnF�� R�"O-�3�Qv�8P��ڪC�b���"O����iŔ�� ��� <���)�"OT���[<��l�W�$6�bT"Or�A����\YU׆:���v"OT����Y��V��utxC"O��E�.��%�J�s��4�t"O�M�HQ�s.A(g��;�~x�"O�P���}�h����
HS�i+$"O ����Q�ԭз'�p.��p"O"�CF�!�l�`��r���)2"O�ij1,��bo��@����Y "ON1JĠ1V,f�3b�X	StfI�"OVx����^�ɹ�q��b"O�`���4	���b�F'�t 0C"Ov�5�_��`���(EtX��"OB����~z�c$�6f6@��y¡��C��qb-��|"��Ю�y��
�t��c(���x���X��y2�Ұ�\Y�D<cB�AR�@ �y��@J�9��!αT�J��v	��yr��f� y��F=H1��5ƃ-�y�Ł1� �k�gսB��dK¦���yR���d���CІ�:W���@��4�yR��m�%9�m��9��]{�KZ��y2!��nH����63�2��k���y��C�Ͷ�z�oϨz�>�a �F2�y��!}�85�u�� �U;�$���yr�0.� Q�ACX
��y��D���yb� O�6pc"��{��ꇌ�yR���7:����K�n���#u/���y
� ~������BQ�ݩ#o�X3"O�|� �	3��X��%
_��yq"O�̡V�ȵg�R��kOL��q[D"O�ݢ��G�S��}ٶ�S�D�~P�&"O*�8� m�Z!6�ʇg�6�2"O
�ś W�ft���U'�y�"O�	�d�'�}Q���9A�,3q"O��һF���2c߂1�؄�"O��T��K���R��q�8 ��� D� ���Pi�r0�
�I?|��?D�d�I�;gxFi��g^%� ��`=D��!�ȃof�Ч��8�ذ.0��0<ic"�sH��S�ѣU�@���_v�<�`I�:+_\�AN��	�ą��$O��1s
�'�.���J�T�4�y"e�'BQ����'���(�E]M��`Z��!��Ԇȓm�le3i�.2JA��"��y���̙2�T��ݱ��ɖCE.ЇȓN�4�Rdj��?
��Y�Gbfe��M=bQ�����}D��{�/��O�^��e�f�@��53���FaE96��'7a~!� ,�4��W�D�H�R�"ȥ�y���`���a(і�H�ۦ땔��	[X�`zL){��@����@����6D��;a��0�Yqi��Y�}�3D���a/! v�Pf�6c�,밁&�O��hCHȂ+_p��8Q����t����󖃛!+�n��Q � �Y�ȓh#H1)��	�W�KB�(���r3D�b��@9\���q�
&3�.���:D�T�� �8۠�)�cI
3�� /D�tBQ �:��t��zCv�Cg@,D����GkUH0z�ϐI �xƋ4D�\��b�c���&�
~�4�(��?D�����Z#c�0X�A�	$=���!�)ғ�p<!G ��`#�5��Es[4 ��CL�<�K�-^;�t��ƃ�T�f�Q��]ȟĄ�QIj�b��<3<���`Ԍ����M���	�9��rUfP��>�ȓY,��D�v��i�s��I���Pj%��
A=��A@@ C��y�ȓ7�n��bBN~�x1�ҏP�\� ܇ȓ'��[�W�=��3q@Q��ȓ�F��'�P�z�R��Ȋ�di�ȓ0��9�j	�8�t1�U� �f�ta�ȓy�PТSB\�քab�ơ�F�<� )Z�Ii�0���>Xw��*DKNm�<�Rg��/J-*Rb�d��F�Jb�<!T�-"C9Pf�,z� ���z�<!l+�z�`�J��g�p�����t�<�E�֜8�\ɳ(Ș 3�8h
t?YR�)�'Z<���A�=)�$"�T�E�X����ȅ2��? 4E�1^	��Z�b�(eG2n>D0����;<xM��+~\S�"ȡO����{*�Y��J����]�D/����c��@/����emܸ�c���"�����E.8���n��U1������f�u!�`�ȓo���ğ�"6z���+C�q�ȓ|)\�Zb��2!4��s��)T ^h��!���҇��&�0@�X�Di^чȓ!�DY�㌛�N��#p,J&����v�̴����U��Q�!Ϲ(����ȓ1)�Hb��4�t�J���M��ч�S�? �2p��T�Hu�f��g�fyh�"OL�siӉE<�xz�iƳ}�h�؁���A���'r#�aa`���(�,�5Z u��T��wK�Q����9�u�����!`�\���Op ��O��b�(���I^ ��%�*�O��ˮO��k4�$!� �D�e�	q�"Od����)�p�
�D-	���
I�?�¦��m<���D'm�^��b�:D���,��	 �T�(<B@9�Ɔ�>Q���ӓhqv�u!v��YQL!c C�I X��EB/52���҅�6M��'d����Ϙ' h���[1`Dɕ%W#"_�ī�'Q����*	�-h�SE�Uv"2�{��i��yr�A�p`}�w@M
>��]�,
��y�~�8RӣI;z�� UD��y��73��Q1TD�C4�)���_�p<)���R (N�j4��#>�xPI@� �!���VN�j���h��u(厜�v�!�F7~��\[ �#U�.��'��W!��wH�R�ӭ!�pa��ct!�_�v��%�fH�!k�4�B�/eZ!��)!�\����W����N�(Z!��9@i؄8VɃ33��Yrsn�&
�!���.��� �雂l�F=��-�'`�!�D�!m�8���B��H�s�Mάt�!�w�v٩�`��v�q)��ǹ�!� ��${fƍ/n��p��=A�!�Ĝ�a�����-�DXH���)�!�Ė*g�p�P�ôS�|�A�F��c;!�$��`��=n
�{'6����/�B�I,V��Ren������A��;R�C�ɩTBU !@[�kj���V�P� NC�+Q\f|"��%���R�h��nL�C�	+���@�dжnXcb�P�W4~C�	$G���aL�7?�d�_���g"O�ܠD�];����� ��T5�"OX!��#ρzvn��`"�/
� @"OL�1�#U�`k4B�=)����"O(���Nz���&�5&�Qd"OD�YbB*&8K�<=(
�"O\iZC�ea��c�k�,8�=�"O��"N��:Y`����%E���1"O(@�h
1p�i	<hY�%"O����Q�X"���f�	(����V"O�X�@���y���.�:��H"O�1'�ȈE"�M�*m���4"OzA�E��#,�\l@�,9xh�X�"O1���1b�*���J�8L��7"O
}�C=�1���C.GT"+�"O�|Ѐ��4$�F}��l�#N綝��"O��R��7_D)�k�m� ���"Or�r)��s�s�J�!�uX�"OB��O�M#@$cFJX6|��p"O�$(��6>��F�D+b֎T�'"O9S@����X��s�Ͳ%b��h�"O�}2gϖ�<{�!c��?8G��SD"O�Q�#�}�a�"۝><8�"O�q3��!?o:��V�����"O8`��⌎&�B��%�
2~�X�y�"O�%tŁ��e�]*�6���"OP�1��6X�2����, `!e"O����o��M�4)(�@ӡcXI�s"OT`��S�(���# �
��1"O�$�&D��tL�����xOF���"O� �}Q�CS1I�b�@�(͟4�X�3"OP`1�)��rZpY�Un_�^��	�"O��31JmZ�A�D�V/l�`"O�٠��{�搉q{8ͱS"OB\��˝�D���t_5"O���+�a��d�*�=Q
4�4"O�p2�Cߔ8��CpjK�G2��z�"O~�!rM��jd�m��.h��B�"O��Q�M˯#�><I��-�%"Ot��C˗`k�A���W�Z�%"O��2�&�1�D�DEn�(0"O� p� Z�2�H�N$�ι�"Oڈ���-(�phFC�]*��"O,�Ң��5i�68�t�X!XsR���"OĴR!m+$�DՂ��p48���"O0�!�F�P�� ��� ����"O��!��/�>�z����s�C�y��(bbF�f��;r�̃��V��y��>cdT�ߪ#� ���y�ˆ4�[rဈ!k�\�����y�0*�����MقI+2�����yR��}� ��UL�:e����,)�y� i0^��d-J:/J�4`UM�&�yb刦|�J��u�O���}���\=�y�Ǆ�~TJ�B�g���5���y��P�PVUd�R?a�V�8��	�y���c<R���b�/l�y�4����y���JTQ��lF�7��������y�H�%ծi��F�A�<�k3B��y⋍�BJ$2�aN�K��t��(�y2
S�#��+���@�� �MS��y��A3h
�a�iѶк��I7�yb�R�xYM�UR*��@���yb��>c���A*�D�X�B˕��y�-�W|N$"�0>�Pc�撳�yB���23$4f��!�W7�y�G@9Vݡ��77�E�b�P�yRbA�B�mp��D<��u�ح�y��F*o)��
��䃢 �yi�U�hZF,_5I���4c���y��]��D\X�B�
���r���y�N��p��iʆK���%�B�� �y�EJ,M8�h��L:���S�fH��y��_r��C�#���(r�L��y�ʒ�-)l$� _'B����l�yR�L�gc�ԓ�jڋ+�`*����y� �m�\ub��ґ(���@ǭ�:�y���F�5��]&��7�Ҡ�yb)�"�pb�#(4�+�S9�y���Q�(��oīX�MHR� ��y���L}�u�*W�?��q��'�y�D�l̾�"mi�b9�0K<�yB�ڂzfp0"_�$� V)�y��?�|a§,!,H�Q�I��y�lԧ��MA�F_�cC�c���y�K�-�~��ì�Wބ�1�!R��yRT����AX$Vz�$��g�y"�&L��Rm�6G��1P�I��y�	�)P(�Y��ǯ3�r@õ@��y�*K�l���kX�'-2��d���<q�����V�="T��1��R��!�I�|����Ã�!q&D A*�=d1O�D���!jP�S��D�}�"ԙ2��r<!�ٕ �9)�_�l����@� 2,��� ��(��)� ���$�7��u�
�RQ�l�@"O�����@���FD�yL�q�"O@����Ն��0
Y� �����'�n���'�&!@�Cߝ6}�	P%��Y(�9��'7|��G(͍N����H�R#`���'��q�AЄ=�ȗ��H��e��'bbm�q6�V��&N�>̝�'�t�Fy�����S�9����9D@�����b�!�d�W�����ۈ4  5ɧ�Q�~��	q���gHK��MYu!��C�Hɚ��2D����`ߤX�L$��#� W"�u-,D��	��3��a�K�D�)D�X	�bbJ!s�͉�Jp��'":D�0�$.�
j���r��	$�l�Wθ>���d��-hd��>8Q�-ɔb��}<��ȓfA��ݪIb�x�d��r��An_(<9\h �����@�Yȅ�A�9���~�is̘1gh�*u����b�0�f���%kLT�rH�1V�@�� �
��H<�O?�Ʌ>��%PC �� ePxj��'��B�I�+�@�в:y@� �ȕ�B�C�	tr�A�3&J�B�H�bF�oC����)���8�� U��'�J����{h!�D 4��T�qH�Ⴄa�g!$X!��KOd"�䃑D���Y6`�/D?!�E\$d��W� -V�!9�a�/0�|��x"���^��iH&Z�t�����8�y��.���������A������O`�~jqKE�?�F S- �KR�3e�VI�<qG녨Uy�E�P��l�@FNI}[�8�<1��dπ]��lɕMc��:FGN.-$!򤅘Avh�!�
!o�+&�+B�!�d�^",	ؖ�͌9U���Џ
�Z��{B�ԋe��H�BҸo:%r��/i?�O ���ѱ��L��J�rvn�2�A�?J�!���'D�
�"D�5Hg�ՒB�!Sw!��*8�q��(hK�s�/K$lX!�d�.&�R�p&�N�мh�o�?(��E{ʟ�X�F�(#*ĕ9��Q�|��"OȨ�v��t��ȩ5��>9々���S�����:2Az8�C��=����W�Q0I�!�d$1h�	֋W�2�٠ ��t�$Q��Hs�S���ѣa�Ɓu F�H��ÑfW����:}��Ƴd���Y㖏R#�eh�hѫ��I{X��렮̥7/N��W��2����"D���f)�<"�&1d+θ~~��I%�"D�x����*�>��Lr�$Cw�<D�CǁD�1��8H�A�8l׶H8�d-}b�':19���>M�F�����,m�5`�'���	v��!c0�À�P�'�.t��'D����E/U�xAx�&�E`"�R��F�O�B`��CL�*r��%�Z�O�dA��O���ŏY��f��2�H�
Z�3��x�mpy"���r�ܚ0K�+�y"�!^,J�B�	0;֊5)�bJ:��(f�\,*s�b�`(��'���鱅��+�dl�$�ۊzFNd�	�'�D:�)����L@���~U�K������<�H<��'��n��y�r�\$�B�I�x�9$�Т5ߌɢ���J`XC�Ʌj8�[�jT0~�(���/�5X9B�+2X�k��G4S�8-w&��9���k���� �{�J��L�I����R�"O���q�З��`�g�#!t�@rQ�܆�������Q�G�`�����7v�,������� ��Zć�Ax�DQ#�ۺ 4�݈S�iޡ��L&PG��ņ��"GhP�'b+64ў܅�S>����%�h�b��	�+��C�I62J�YPP�ͪ{�XHBS땝���>ғ^�j�S',H�%��8 c ��#�H-���b�X��L���ݓ$�
�+��I�X�1�4�,�?�v�S/+��)֤�r�05*�t�<����6H�l�diI>x0���JyB�'da|�DJi��[b��auB�gdN��y)�\-�C���/u<����Z��ye[�nI��ēT���b�ƞ�p<a���!c<�+R��y��@�6�:z!�dĹ8sV�!t�&c��af�)P��hO�F��v�Y�a:���%B�L���"On��blA9A&`(6�4z��ݻ�	m�O
 �aĊՖW�0���M�\%��(���yBJʽ�f�8�@X=:�@(�4̎��yb�L2~��`�4@��\�zȈv̘%��'��d%��|Z��ۧ[�ԝ���I�i���QPN D�l�PnR	Tb,�	钨wn�R%%,D����Y��D]>�0ɒ��)qc�������'	�h����< E�����e�~�x�}�7OHc�H�OT�U�*.	l*��F3G����>QN�X�	S��O�2��)��5E��3�R�*c\���D{J~�G�:**���'�ʫ�,P��]�<�Sa� |��L(��&n�X5�'l�N�<�C����ذA�Q�V���IJy���s��(�r����o2���ԇZ'���ib�'t!�d��}��AA��Cj����F�/C%�IR�H�<ѱ�P�\�0Gџ>8���Vk�B�� Y��Od��4O�YƉ�(t^թ�a݈'w|9��3��8*wn�H,��
��nZD�����f���N�`Ю5EFL�1PA��y��%
�p����Ҋ̈9�-���y���:������y���H
�y�썏g���
���&��CR)�y2ꛁ(kd�*�힒�2EZk��y��(P�`չ��^@�.MSbc���y"l3L
8ͱ jN<`h(�	��y2X�P)|5��
P>�0��g�,�y�o� s�u�r�[�J���p��I-�y��=�\���5e�8��h�'�yblJ�d1��꠬�4 S`Rc-��*4�0e�N&d��)��@�SDȠ��$D���T�4E�I�+M	���T#$D�����˫Dx:dzjo;r��&!D�p���ɸT^��#��5�^ԓ�m?D��J�J<)������'2��`=D���Q6w��9��/�"���s�=D��ꇌJ����q�Js�5��I<D�L!#��#���p@�\?-�ܨe�&D��:1g��p� D����'>��v"#D�T�G�5sߴm�v�3x�P4���"D���tlM�|��X�!أ;Z8�B$%!D�@����7qR�*$o��]l,��% D��(���t�bi�2��1&<���+D�|����M�]��T�@�̼t�*D��	�FVu�PԊ�f�;2�ƴ��n<D�([�,�r��!
u�5sI�0�PO<D��"��ϊE�iӃ��4�t�;D��[d�T�' }:�Oi���{��9D���#
Z�*GJO$�L���/2D�Df���<9jdx���S���R��3D��4�Z1�(a����	����0D�� �x�3�D�)5t *2"��k�y��"O���f�c��s�@�c88s�"O�tcv��

|������l(.}
�"O�p���V�m �.'-j��"OJ���->0v���MD�BC��*�"OJ�26��	@D���GNW� y��"O��ؐZ�}�6�づ��-â�ӕ"OK˪@LBآ&M?�ʔ)��]��y2f^�_d��80�Uˊ��HF��yR�]JJe��+�+F`�l��5�y(�3�$�+2��E���9�i��yb�]��b�y3M9f�ب����7�y��ލyT��f��4^�JY�⧙5��	>n��.zq�e;dvJ����D[B�НAAZ���Xs됈-k!�D��V���ct�:p���*D2~J!��Д)0��y�I�9'�4�;�

�sO!�وTsޤyT&�*`��p
��U�{�!��u�%jBe]�S��XP��j�!�$�@�-�W�8K`�Z2u�!�6�H ZÄ�(-,�-21	M8N�!�D����K7#ʻ���q�	�(|!��E�S^"����ò&��$�bA�!�ēS�>�xb���y�����d�!��}C�)i�&ע)�&���B�	K!�d�UB�CB��s*f��W5!�d�����bǿTvv�)��E�^D!�$�d׮��ȓ#��42� e'!�D@�e��a���޵Cyp�c�˒}:!�D��u"��s�哞aix�ڕ�ԥ<!�DС|H����݌TCN��BĊ!�$=����%��e:Q#�+!���P�Ό#CB����ʤb�k)!�]e����Uc��p֤0!�R3E>��iK�#X0uc͊~8!�$ijlt)��0g-L@����4�!��ߺ3z��� �4;�\�*#(X�v�!��H�>������S�R�ĠH ��/r!�u�5����>I��1����.T!���L!*�l׎T�Zx�g�N]!�$X	B��]�WNG�&��l{-�P-!�DB�6tP0�7Is��;�̙�!�D�#),H�tMV0hxY� �(W!��Z$�NQ�t�\.Z`] ,ʨ�!�
5k)��Ü�]9�B&�F*�!��P�t�`tR �^{�E2�c�w�!�"R�^��wΟ�WV��A'��c�!�$�'^L�K_3]��5���R3�!��'h��)PA�ֳ�D�RNI�L�!�$T
��#voY�&\4��-���!��D+<�ꔲ��D��D,Z>Jg!�d'WXp�Q�K����7�зm!�E\���!�C���܈s�C�Tu!��F�?�`2&̀�c>N%�%��m!򄘮p���R$�w6�0i�Ȓ�bG!�dI`N0<a�
�*^ր��n_#]4!��*k�:�L˥a�\�xS΀( !�C�wh��E���H�-!򤕆'�(	����(K�*�b��1;�!�dL�$�d	+�"��#���3��v�!��
.qr\���c�c*R웠�\�@�!�dO�Q~�����)Dz�'j�i!�[�C-��K�S.?��:�k�>b\!�D�8�&,0����<bg�)UM!���(n	J�3�H�}[@)""CA�R!�� 8e��-B�hr�Ə3!�D��"O��ς2�V-�f�� �9��"O\�3��y�(���b����"O4�9r��M�`��ޝc���:"O��(� �7��S��Ћ��x�"Od]S��,^Fly���OV~�`"O���3�Y�ɴ�FM�1�L���"OvX�5k�@~���@7.��|�"O���c��1t�4�ܤo�0�"O^�+F.O}R*��)ԲWy�4#E"O�Q#P�4)���.}BQ�'"OիD��mު���G�Z��P"O�Iy2M�`vX��愲P{�<�"Ov8�M�9�@���Ĉ;Z�:��e"OP��D� �<�ScF��*��2"O<�ف�K�U�Z�p��4'�=��"O�I@��N�\P�e���n��q2G"O��C�E�:� �Zc�Жn�$�"�"Of|�'��2&��q(L�Jv����'��|ЖA��T1v�+Y�n���;�'�MZUg/_�2��i�g䤀�'���䛆���`#�Z6��)۴ ��t�P =�O��D��6[{EJ�
���j��'�Z��®j��	5J�r0Xe��%؝÷�N& [�B�I�x�����E=?TpIw� �z>d�]*��y���:a���A�ܼϨ���C�E�
9`�����ӱ��Q "O��`"T>h��:D������!^.N�#ش[���R���:~�&���'i\тj�*0̒�ч�ʘ�dh�N8�q�j��x�̉����4یI[ԭL=BD�y��+]E�{���D��➸�F�	X#^c*����';�n��(G2 �K�k�7ێ���.gp
� b֟�1PB�\Kmf8�3�+;Y�%R՜|"Lê9\�5B��'���3qiF3>�R��FX0$���C�'�l(��3Jj�rύ<Q�����_.���N-#��ʏ>�ڥ!�=���"b�'����c��T���� -���A�)*^7��P�ŝ,�1�Ҋ��u
֍Ef:<:�Kx���4�QOK#-IJ�����m�Z�t�'��Aje鉏��(��-�AV:�2'ݞUc�@���1>�6�D��-��q�>�Ah�'��O�έ#��\�7��D���OA���h��Ҹv� �{q&О�@��r�X�� �;�������q�˰lR�O	�P�bf�X&����'����W�΍ gR���E_�3(�0s�'���8��_\��YC�ȲE�Q>9[�o�zE��r����d9v��Ù�-�	C������ۘf�^H������2e��J���Y�e�XQP)#W�����J���B^D�J��1��:UbA�yl�SƄ�>���DQ c:��������jR��C�x����^+��l�1j@�$����/��~�'��P~1�}nZ:��x��_rN�cďP֢>�`kL���gAD�(3D�nNP��gF�_��OM>���3(�4���@0}<x��I.O4i�wlOA*��/ l��Ӏ�'���	��O)n�
,ضOѽh1� (��n>a�W,SHX(+&�@8{�f�5�O!caF�8�']��낣R�y�@D��O+j�|���e]�� �'kD�D𠊆�G.W�ɫ�#�p�Dێ_>�Nؚ.ծ bí�5'�ZF�U�u#a}��Z��Jc�EZ>wD��8����M��D"�۽%/~�kg4����>��.�d��>�I)��)��*�0���p��-�>�<��C�+��	�c*�����P�9r�؇W���@w��| �OS�<i%K�[��I7�.\O��֡�;klY�$�Q�xA�aP؀3��J�� �/ǐ%�1��� %�"���֡Ժ����ː�J�����b�!�dY�֜�!M�+������WĚ�A��׈1�riK�{:l�
�,حޒ�I��Hujx��I�ٯ�~���"v���6�O����4���il�1-�F��#�Q��Ё�I�dZ�9��O�/89��M��c6�_�\w~ '?�	�s��� - PiPE���߁��"<1�b�g�	�'��ƀ���?��	ѼY����K�rf5z"�_6u!��rX豰�1lOf�8b�D�F�\��B�$�a'H�	�@5"�!R"tUQ�g��q��� ��G:C^E̓:`����jX�} �`k�-��1���	�mk(��V�Ov�A�<�̈-�8vI�`��6��3�/��T۪�Á�V6	n�;�4B�S@����� ���?)0�ٜ5m�x#�O���� �?d�8����2O������qt�Q�_f��eis�۹����� ��k�Bڝ!j�!�A�4L�����<U,��1���<96~�J���IwfLKr��Sr�tϻH���a�\�1�6���-G�&�a��]7��+D��0�T�9��C��U��?sNT��f4d�q���#�o �֘b!�$�I���iA���9&�Xu`D8R����d����h�jӵ�?IpΙ�2HnHAfN���asMD�䘭(��Ff������5�H��g�'�L!i�NY�FH�Dc��9>��Tk�}R.O�-لtb�{��ܟIW�)��Zl4y	�,��h�:�#ǈK�����擖b΀��䖄$l����N��́����3`a��Bט{8�O����0�p����Q91B�`�� K�#K܈�2���$Ւ-�s�!D���2���`rȡgjɟ]�NE���Oj�FG�+p����թ��y�dx܉R�I_��i)Re[EeN�4��6#B�O7p4�ۓ"�l\��	�D�P�䉶-Fn���קnwf�x������ڻ_�����A4�H�lt�_R�@����ϕ�h��� ?�I����b��	� :�w|�0���M�\��T�h���\
�-#$�,q A嶭YG��3
�Vs�b4D�|R�Kj$9Q4�[Z�s�Q��AH<HԆ���թ5���,(D��8戅#"������s�2�Koc��X�����t�yR.�}+�mD�ܴ��6o�$�*E	"��sِ��ȓ;7���U�<3Ǧ�:�*�
�d��3�N���#3�J.Q�V� �k���@�b�p����C���5�ҡ�73�}��456� �H�9��5���	e I[2��p.\�}ז���']�s �UsP�c��Ta��`���$�,G�%(��	8+И:�ꎱ��)�%P=��@�wd����[�B!���_βaq�J�w��Ā�BF3q��Kٷ'&:uR�W��L�8V�a��M!�/W�ʰ�A�Y��e@�`r�<�Ń�<��(׎l��,`6ᗪ[4r]�,�s�`!��NL�ef���×��hOR����	..}уc�����'*m9D��a��� ���g�pA)���vz������&	\�藖T#p`Y�G8�O������R����dX�;�䉊՝x�É�Ep�+ek��S�B)��J�<57�$+G|�d��>Р'�X�v�x�{�H��y".�:C/�貕�_�5����a@&�Ɓs��,^��s�.� 2��W �ͻ_�H���\���($ih��`��C����0*AB���F@�(Żc���79ò�D�f�9.R=9�)�g�h�j]9��ޜ6Wę�`̉�Yi(����<:g��S�A�6��D:Q�U�U
�(V'$���!��\�&tJe ��A�`��dW$\��&�		lR���D�8��'Ҹ�3��,}�£�KP��U�2P��.�TQ+ H�l� ��c�<Y�!A�RaI"���w�~�pȟ�D!qk�<���#z����'�E��8%��@�e��93�B�'�D-��͐-R�s�&W:���"l��+���P�Q96j�|"��$�p�06h4@Y,�r�	R��<9�D�B\&�R�)�>9�(;2�l���}�������F�<�G�T~��R�#J<e2��OI|̓<g6���<��:��Q�O��NQ�&�&���""OP�s&�̼/x,"�ՍF��г"O�����N&N&�J�CٴSy�=�g"O$��3�#���c���=���)1"O�$���Z�Q��_wa����"Odp�cf�+t,Y���.R�0��"O� �0)�	V%z�9��w��-
�"O��bU��4Dr�E�*O�3��b�"O�\�W�F�1HV,� j�c�:�;�"OT�u L���8��i�7r�n a�"Oj�q�㓋P��2�hF�~�XH�0"O���1NK�1��i��ܵ,)b� #"O��i`*�P��}Iw,ۖ��5S�"O�(�IȐ�R��ԩװ&���6"Oz�{c�-=qt	qwG�7e��Q:�"O��1T,�&X����dĐ"��ik�"ON�J���?��u��DG���z!"O��3���>o�$�atA�9kv��s"OHuH��#q�TS`��,�Q��"O.�K�K����mZPa.��e*O����-o.,cS�@�!�D
��� R�2A��1�x�QED�fK$�[w"Ol �_! �24���*�e"O�A�wҦ����U�/٘��t"O�!Ļ
�8�KdP+w��D��"O>�Hpo�6�,E�C-<,��"Oe�ƆA=���!��p""O~�c�k|Th��@71�ν	"O�Ƞ��B;j��f��^�Vݨ�"OjPjU���4���͎hҰ�3b"O�dQ ��N��ɒ���MY:
!�d��i�e��E�"��+Μ6�!��-{�j�"�Ѐ(��ܘ�eY�8�!�Xt���GMe�����d�#�!�d�� �8yŏ�4^��1�5J?!��.k4RŚvaY�V>��Zb��		�!�M+J�&bѶO2mY�,i!�6d���aH�#$)���P�BR!�S�]����F�#��"'9[y!��0U��H�3DO�j?�1¤ܤVM!�$T�9\�ID�6��Œ#"!�D_�U�����q�i��cρm!�D^�$2��ajI�|�20s���
>!��
eE���� �'.BT�;�!�П'����B�L�<0���ف}�!�D��DV����ʖ&�����[�!�d�)R����L�M��UڀoO5�!�$ֹv��#Y-��UR��5!�����lzF.O�bl�1��{!!�J$y�l�1i"�%��. ���'��Hå�kL�E�Έ��#�'I��❳aDX�Y ����'��,
W	�zpA��K$��b
�'�t���ɓ�B�4��씈��|8	�'���a�
!X
,܃�iA)Jdy�'�Py����kF��bMO,~E4���'�Y�b��5O5JePRb��r�ڽa�'TL�ǩV��J�A�M�������'7h1�(��n�P.��%;���	�'Q���!ώ�7��D��M���B	�'Y� ��Fp�,��Ƌ		)jB���'F��ȣ���O��Q�	؝y���'y����P��G ������'�X� ,��o|ݘ��\Rl<��
�'����C�.РR����eP
�'��Y�skۜR��]�eO¨v���	�'U��f.��$�P��i�\���q	�'�R1)�d &�����/B�E����'�ei�/N&wU\P)'�I�4�|;�'�ʘCC	M�)U��9`��*�,T�	�'�>��l̆{�>9���# �n({	�'=��0Dֱ/t�K�$�����	�'(F��"dƊ˚��v��
#��q��'ݜ�cR�2ź<*A�� �j�A�'�����'fu`hQ`S�i��b�'���m)w%�(���@�y�(��'�.m���Y&J`[�WAE(��q�'s�*ad�Y�����t� �[	�'�D�Ã��
�����s��d��'\�(V��G>@�d�ib�\��'�`�@dꈃR\ ��AÇ|���'��PQ�K!�b�K$DۻX�B���'�e9���2:�I���X��8�'�^;�5tH`���C�_�,��
�'I���"C#l������8;"�

��� d(ˣ����SBA&/���0"O�҆͗�w#��3�ЂO�l�*e"O��*$���*@��-�@���"O�i���-�����5�D�X�"O�@Yta�6'�92�K�X�d�PD"O��2�I/��I�#CB��@�"O֕��j|=�Ba�;qb���"O�9��L�1��9b��6Gb���"O4�p¥�D���Ǜ�wY��"O�9u�_9ŨU��uW�%��"O�ā�TӶ0�����MP��"O�x(f�2BLP����V_>Ԃ�"O�옗�R�b����Ɋ&>�u��"O�}AB�A���C�iL0�,�*�"O��@s�Cc��e�a�j]pD"OBdY��-[���X�h�8wC�9��"OѸ$�
���M(	+f�`p"O�a�Ƒ:g�$�Ad�.�%e!�D���
Gf�H�9F�1!�MV<2}�Ri�5��|i����q�!�$���1� �����Q$d�?�!��(,�:Ca�H/�D	�Ă,G�!��1o��}��Z�l�3A�!�
���ࢳ$G���3!�3QV!�7?�<�6՚`���Ǣ'?W!�D�v��\c� =e��]	��Y,8,��n�j����I7����D�?�웳OW
-�d���Ϲ����b�>-�I�V�@�K�zm��ҁ�h�< LL�U�<�+�-r�4�G�^`}�Iߙm����SdA�A� 6�S0 @�2 �?if��M���
C�	,k�" ��$��lRp�s!�9u����V*��IO��
�u+a1�.�P��$�E���R/W�ऺd�_4a~�o�
��4�`�@j�i���E���W�;mc ��!��H�QI�g�ܓ$ͬ�>�Ґ��\�˧/9��!6�Z>�6K �q���Q���?a���>�.	��H�@`�B��;�Ob�b�g[:��d�y���-zd+��ʔ�Xl��0O��!"F���T�'�]H����tˁ	W�R #"�P�M� hˮ[\jIQ� 1'6����e�8�����+�@�X�n�V�R F��;..>�KU	�B})�hd�1����Jp��ru�>��oi�P����"~U���>-�>���	�Q�M+Sǃ%Z	�Bgߡ@��L�d�]�x>�E�U�
$q�Jt��7LA�]�O��4h1'�0IP`F��H��@��.��#>���$ �H��i�.��U?Q��j�-2,s��ݬ3��=��+�u���:Zm45Fu�3���_��"���ʗ��
��ɻ!Gp�h!��y�!�Ў[�O踥��)@0_�8Li�FL�f���	�cV� ?[��*CT��К��xN�0g��HZ�;�ω�'`XΓs�r�Y�$�'�����	P㝼|��s7�օxpf�
��FS<�mSV؟h��.X�B�ܴ0��TjV�./���A+��U#����fa��ꀂA������EV =#��ܴ9I^��QɄ�$M$ ؅�?HF���ɹ%I.4���U~BI�� 9��X�q�������~�E�|è�#���6\\i��ɿa�񘅧\������h��c���5�[i��Ohd#rW5}�6�[!��3d�d��k�<w��t+ѵ�<B��3g6|p��D<c���#ׄ7x�#<����*l�LȠ$-ʧ^�T���f��Y���Y� �� h����e�Nw.�؃�Q*�����ً^U^H�$�2}��9O^A�&�K�ܰz���Ȍ��"Or+��%<��A�.h`x`2�6O��"�B	J����u`�Ƒ��`GK�ȎE��X��� �lK�u�:��!&?F��[�m�#�h�!�*D�Ԫk�	�*�MB0�pC%:�o̬d��g���$�|���R�6ej���)���e��x�<��RHR˕=ڜ"f'�N�ZT8���"ǲҧ����ޥd�����_Ԋa�I�"fe!�dǅvm��	���8k�t��U��|Z��͠��M;��7lO�YR��U!%����n� .q:f�'?T�T���� T-8���4�~��Տ�.1�����'�r����D?���QkX�M�A#n�<�RIŷL��\�ʀ�H�Y��ĉB��K5�,y0%
��І�Q9Y���h*�rx��
a"O����H�M)J-�b���V��8��?:����4}b�=�g}�K�5N�z%y��9�ĳ��V��y�/���آ���?�4- �����M���]_�<���=���^� 4��{� �kc�=��[/B;�� A�ܰ=��G�,ph;���O��i`䅜^���',N�Z�]��s .~�`<��	��ڱ)�DV�&���È�C�Jb�8�p��$(:B�>i�N�L"FD8�.ޟ%��i�4�ڿ��`���-�C�I�Y<�Y�t*-o�x����>
���c��K�X�&� ���F?N�B�$�L#�w6�����U�=:�k�un܌�
�'G�C�؉�2��0L ������dʄ�x�j/�ēc̚!k1�T�]��ON��@5\ ZC"[${/RI��'jLp��� �����$
ΕأB�c�K���0qB7S� � ���18��'F$A���G�;�l]  �_k7�<+�r��e �X�T�xrf� �R(�t)�SJp3��)ﰅ·cY�vI�h�ƓE�q���9cMv=۷�D\�8Q�`�7y�B�O(it`�5}�L�#N~λ7��4T�R���Z�*Hr:x�ȓ��a����4q4ώ�G��l5-�>|z� A�'���a�H��ȟ��$.7��Q$ߦ�r�E�_
�y"��-K���Ƞ�%�5ru��1�2Ѻ�XFDJ���#V5��1+�Q��IC�"Z�|�qlO9k�����>�O�ʱ@�6P�BC�T\�@|��،xQp����/7c@	�H�Wx�!p���^�c�	Y�p����Q�?�R���g�K)��$lM:LI��'cǚp�Q��$v�� #�� ��ȓ/Y�Yt�	�I(iq �����oZ3I���a�')	���!4c]Q?7mAt~���ي#���a�ÒF�!�d33܉�E�F��C D�l�@�Za�����3
�!�L�31أ=a&F�'��ix4��>+r��H���nx�lhtc��)w��p5-0nzl�"� �Q��1:��T�8\�q�@b
&(h�x%K_���>]��z3�C�<^ͳB�"�Ȑ&�(�7EҖGp�Ŋ<Vc>M���J�|\8ia�Q>%1����A�x1k3�$LH���R<D�D#d����ؓf��xu�L�p��6G��1A�)?<kvP�g��x�A�}�C�چ>����Rq���V��q�D¹?���"	�'��x8��®S��[���?pY�\����D�6�Z�J �F�P�;�ŋ�iVdhH#�c� ��aɖ�.����V���	�?�m@�!�*3�L	0S%Z��X�o�'I_8��#d_����Iq	ށ�y��I�{״�:�GY�A��<`��޾<\tOL�A`��{u��r$�[�� �����N�~��%O6)�0S���y"'�>hf9@F��#�l@@��Kx�����Cy���y�:c?On�;�Ȟ:Y��{�$ءT�F�X�O��e�Ń$n"�ҖIN	T��r�G�R�R p��¬o������7�hs�cF2d=�U��DR�Fx�y�#F�f8�A��q}�o����1P��R���p���y�!��u��b`��)j���G ��'k���gN� 0�?IS�� �����FÆN`m)rk'D��A7F��&�l�����1\=��+8D����I'Jl�]��ŀ< (Y�G:D��ە%֝RK�eS��$�<%���8D�4s�o]�] ��9��J�%�
%�R 7D�(��e#w�T�CPAɍY���� D��ӤW�i\�I瀄=	+.P�Q�-D�P���(WW�Lꄊ��,b�0�wI4D��S�ހTSj � �E�D)�Q�?D�|xehCm�2�sm`�u��9D���bK�* <�C�+��z߰iX��0D���Q�.<�a�#`E"��0�,D���w�#"�Ҭ�'`_]<���O+D����$[�Q��8������(D��i�`\�#2���X��'D�4��g	�Z�
	��#��X�neZ@n0D�P.�+(����E�T�R�P�,+D�� ��0�s.��Z6K۹"���#�"O�x��*ȳu�(,˷��=�(\�"O>H�  �Z��P��?��ĸ�"O�h0G�/y.�p��L��R�F�cF"O�G�*2�@i�kѨ@q���<�ū�b醜�I��Z\juo�u�<�1E�3pH�'EJ
C�da*�Mz�<�4(T/A&x�RqI)	!.~��B�	>I�<�ӆ�'&!~�Z���z\�C�I=?���Rh@�z�
�C%ɿj7RB�	�j�>��w��2���SP���m
:B�	< cN&N٢yD�����*<<�C�(#x����U
� ���N��C�ɧ���@À&$�.9��NaC�	,~�H��B�.,:��6*�71��B�
,<N�s�
�n����dΎ:q�B�	�:!���6H�֐�T�R�t��C�	�q��[��>1�X�b�Q�[L
C䉅14���dM�O��+�䌆(&�B��M�ZD�g+ \���E�%LG�B�I�U��i b��G��y���I���'�|Y����{�P�QA*]�jZ0ʈ�͋�p��iñ�<�t�`�O
�yR��3���A����
6�$OO��yR$��D�������t�ʭ�딟�y��,-�X�����|��;���yr�P�f����aa5o��a�r`׋�yBe_=�r�2��I)anjP�5c
��M��aQ����ȟ����P�P@��J��(ĊJ��9��'��𩈼^Y���%��D��l��GW��+��$���]%?�JR՟�������\��͈��c)g������͔��� �3���r
�'��=a&�<�> �B��1�c�O,m D�(,)j��'k�|���"M�li��oԓ(R����Iy�%�ö}��T�h����F�Z(Q��!�F Ŋ�����N=l ��2�k�k Z�S�O���)'@G<(9�l�96��,���p|d��lyb�O�~1��5#l馅�BZ���h���	 ��0J�O�Y8�ųVZ<�EMX�7�Ȅj��<� �4cyֈS*1}��Tɍ Ma��Ԍ�#\H( c᙮�~���dp�� �|��ɒ��pJA�V���[�GP�	c$���4L-�@b��t���u��b�'ԸO��	����j��&V�1H�������rͨ1��,)jj;�dK�����S��]1�(0˝�Tr�b�J����UcJ� ��ij���*4�l�����\�%��phD�y�K�Zs�<[��f��Dt"�=bE0�u�̲'�&�|z��8�8QꄪŶL2�����s�i#B�pu�>�����D͑_�v	��H�H�ޡX`��!�䝇\��KE�W:���Ui�4o�!�d޾p͘t��;z����� �m!�DԨ}�X��& ��>�ى3���tQ!�R��Uʔ�G�đ��	��O"!��Ȅ ��8�S뇃mu�x�DC�x!��{b��g�^!̰�2�A7O�!��(L�DP�v�O=N<�ؙ% !�$��Wn$�d"��r[��4�ɥd]!�$F�@5��d�_�hcV�a�R7�!�dB+z�D���H	D�	�q熆^�!�D�-"�|��EX[1�Ͳ�F[�d�!�䗸<�R���䊛Y+P���O�3�!���YE�4(Ц�v*|���U@�!��`b���a��"k~�����>!�$�d�y7"�V��q�� ;!�$�-P�a�T�jL4��'n��`Y!�d �TH,3�6l��rBf�"l!�D9����G2z�� Zp�5nbB�I�3q
����/M���!_83JB�ɡC(^��U.L�6����p��h�HB�	�b3��0 ��y�GB�B�)� �ܣU��~�٣�,�����z"O8�bvH�P�4�q2
_�y���y�"O�����ުLՌ�G�#G�L�w"O�beߘ^d�L�7fY�\xԝ��"O�C�
e�J��'��(9Е�v"Ob��F�D�0�u�r'���Ai�"O8��&����l\�@�Hc�3D����
�-J���D���,�[&�.D� �����M�j�+��,~��2�,!D�(�tC�	"��0%(�0htX��>D��hv�͌wW� �%�̓K��`[$>D�4xS U�>�t��*��u�W+L�!�$?D�F'���qE����"O>����;A�qG�Y�|?��+�"Of��Z8�	g`�8<�f�C��T _�!��4:W0�r�'�%�V�BC��h!�X��A�o�!4�0�*�D��;]!��@�08���������kL!�ۜU�~�b֌v�.���_F!��OcU$!J��΅��`#���	9�!��R S,� �u�;H�:�����T�!��n�8Qv�� �h�x�mX%]�!�$]�9v@�%��;~@�'bT�N�!��,;K��� ~ ��y��G�;!��߭oј�:�卙Y�"`�d��%y`!򄐜�$,Iu�_2e��ɫ�˕-T!���,G���.I5=��!�p�J5%7!��<0g&<!��)�(�!��!򤌪���둌p�
�3�
f�!��<n�<��M	_ؘ��%�	**!�J"zP5��-J�B䀙�e�`%!�dS_\�hvǞE3�����m
!�C#a@�}�T)L-P���0M�=X!�L�C�Ȩ��O�2.�H��&��GW!�D�$�֜;�#T�W
�6&�EH!��×|������ 'ؙJ�H�7B!��N6{��ː��n����p�ʣ#!��G���%F©Mj��cD/'h!�D}�T�u)ѥV<�P!�H�{(!��46bk��нkB~Ŋecs!���.Bh�4� #;4�\���C!�$P+>:�5��@�o,���/\2%!���z��hT�/ �\��ڭkl!�DP[�Vq{�Gi�-B1�

=�!�$�|����"���8ն�C��!�,x��+b,�D�0�02
V^�!��R�FȰb�7!�`�+�h��!��1'ʄ(9�GD6]��X-_~xMr�'�! ��D�d�Y�/��dE��'��d�\,w0�M�9��h�'�Ht2g�6٨`�2����p��'V��b!M7��H��,B�C���C�'�v�
Vn��r������m�̳�',d��`"��
�m@�,�I)�'��B6�A�n��A�%	Z�"6���':� wI̿;İ��i��"���p�'�$���o����\��넿E}��	�'�^��V�!wԬZ�`�<uDԹ��':�C��]!g@��`e��mX��'�~�ЖA�7*�p5�H yA��'�
�xC�:Q�Z��s�̌8`�����Ѡchr�:+׌x����V]�<顋KF\�MaA�X�P^]��_�<��J�W���Fo4g���1�HV]�<� �Z0�Q�s�]��E�7u��x�"O����ui�IbgE�k�B�8�"O:�f�0'�1Ä��V�`�q"O�#sᙇUr�@g�T?8��"O�)��ϑg~�)����#̵�"OtyP)�5
.�3���. !p�p�"O"l�l�H� �b
�o��� 6"OY[�MG�6�����O:t��p7"O��#�s�䭂N�* j`�"OdqHF��2��h۷.��#���C"O��C� O�~=����#�-�6�a6"O�(���I'x:9���@�h�|�x�"O���qS�A�:l��D���<��"Ot4-�J!0#d���2I�U��+�yB/B�fV�t���QW80�����yb�["� �����g��d�A��y¡�V^jeK� O�" z�ػ�y �.���@�W0$�c�mȆ�yb�I�,Y)�D��(�Z�mO�y�&TwZ2�KC�J�4$*!� !�yb�ۏBę�s��;�2�A�1�y���gqz@Ybeҟ?k<i��"���yH�"h�P�M��0v~�3J��y�%Uj���R�/e������$�y(�-a��b���'�(E��@��y2#C�^	΅" I����%A+�y�ج��m�di�5�|,�b̏�yR�ԚCD������t�¤�
�y򂘓-��`�{P��@��<�y2��Gv(Ӑ��q��	��N�&�y���J�ѫ�I@�g�ő�E@�y2��ÖD�$K�mC��`#��y2A�W���zd�.p^hHA	���y�R��0e	�D�tԐ��A��yjO�f�&9Atd��h��#�AΤ�y�F�V�
0��.4g%J)�G�:�ybl� �ʡ��
�fiJ�ж)H��y��S)< ]JD��Q$��b�B��yb�ՃI�����j�䁨%F�8�y��Rl�]�A� 7�X�IN��y���$?�!
�ǵ^�6�k�Ꞩ�y�
�+#f0��S<��0��(�y� ܂,��#�ӀO��Ly��K��yb����l���w� u)e�J��y�	Y3BǊT�#!u�TP�c���yҥ`Sу�"��~��x1�% !��/8ޜC����&�p�:n�R!�F&^ޚi�̉=&��IRkE/e�!��B�?��KtlF>�й�4�ɉq�!�do'����V<�(ZQ�N3�!�dߡ2H8�+ь�h��;u<(*!�Ҟd�vpd��6@g�����)!��5J�ƨq2;b���,ˇ)#!�$�0_�$Y��B_^�0��L!�DY5B�α؂��pb9�%�ss!�υ�����SU\��ꖈL�!��*�PS�A�� 	QI^�e�!�DR�Ą[��	�6ᬌc�.ٕRk!�F�u�<��"�Z.��{���+\!� cgN5RCʕ�S�����&X!���p��M�2� ;�4���g˜k!�D�M^�)c�-����va�&c!�R)&�P
ڡ{�I� JgD!�D܅rD������,��g�>d!�� `��D��]����ulD�d�VYS"O� �d���:(8Bn��sq�|)6"O
�����0��u@�/�&ѠB"O�x����.KaDIi +�,��"Oze��'S�,�~H���-q�N��g"Op���hĢ!<4A0D

�&(p�"O� *�h�:/H�{�c��6�`��C"O�� �Z�e�쥃�k�V5ܕe"O�p�V�� :��d1X�bUz�"Ov�!ɔ]*���Ҷ]�9x"Oi�($?}$q�uP�p�:��E"Op�¥��gMTIC3����r"O� P$ɬ�T�&E��.��(�A"On��d]C��lp���G��]�F"O�)�ú.P��J9��5"�"Ox�$ܚm���聪�y��HA�"OZ�9����6�l��ө�0;
�sR"O-�a�P8j�(0�\����rW"O`<@`C=�j�{�DƅsT�t"O���v�C.r>L*�!��@�J,��"OR�Ѓ�J�mS>)�dA��w����"O�|��)U]���(�)	(��p{g"OH�Kuσ>����hJ���u��"O$����G'ʝKC� ��J�"O8�
���$|�3C�+����Q"O8�a�\=C�`�n�
��$� "O�HW�=���P4�T"^�p+s"OKN�m���2��&gY�xǩH�yR��7Fr �pAJ�8\L�dȦ�ͧ�yҬ�R���Y��IN��)K
��y�LрO�5C�K�':7�9�ć-�y2��b!Z� �2)�ZR#��y2�n�y@t�U�2�BR`�2�y�@�7d.�P(����'X���+�yblI�3i��C鄭UH�m�W�P��y�(�"
v����I�!����	�y���1=.�� �|�� �$���yR��$.|N�p5 �)g��p`%E;�yRkâi� ����hk LQS`X8�yR�"rzJu��.�)P Y̈�y���(v]�=U�A�C��9�p%V��y��)e�<� �9-f����Ъ�y"JZ�n=���FKB�1��)k����y��-hBd����+~��`A��"�yr��b����`	�}��`��y� ��z�. ?~���Z��y�	�8Q)&���M^r� <R�����y�㎧H(0�Dr���/�y"D�/`T�z$!�e���YƫI��yR�ۋBX��PA�*d��{5ŕ��'�"%Ӻ\r��l�b�O��xғ٤'�(h���W�Q��+�'�R�'�C��|B�'��OW�q۳�^�0
��W%:a�J\��}�j�: �j�P�k5I�$��%��"��'iB$�	W��?�$�;s�� b���>���� �I���'��I�7u�$l�D�/�4ia� �&v�$M'�0�I�"|��O��YՋ�2`P���'gX���2�'��7��Ox�ĝ�^�b�2��_P���M
B�<Q�B�("z0n�ПЕ'��П������n�,�p0 A!�Kf�'�)? dP��%c�	��La���|�j >m�8���&ܣW�س�6��0�Wo�� �Z#C��I,]��i�<i��W4eC"��wm��fĪ�,Ŕ<r�'�@7��O�����Y�@��g�5m�x�!aU��ukCh��?!��hO񟞸�q��"ޮ��B*�!�T�h��dզ�y�4��O"�T�i���� ��RW�遄�,b �X+�'�v��Mn�����O�$?�4��6�ʙue���.c��|k1�I�F���yE \z�a~rG������hA�2��E/^��M�s��aYR=�����p=� <m��̖�%p(���"�+]���D��<�l���㟘�ݴ�?�(O<�Ķ<��NI|J�Ι#:�<�+\�T�6C��1>[B�y�
o�|}��տ(�c��i�1O`6��Z˓>�<Ă��i{�6�u�|�)�GL� Bp�.3�����O\�O���O~��G�|V�/*@���/�H�E+p���=� �+_c�`!��4'h؈��"^���iϥD�4yU�'�$�a��?!#X?x���`���V�>]���\&"���'���'K�O�O|�mk��݊ ��L뵮�o��Y��G	v�����Bl[YYbn#R�@1F�
�[-�al��M(O6ԃV�Ħ��IL�']Duk�L�L]�e�T�S�S�j���?��"̲!�d��Iϟ%>�҆��%Ơ�e!ϓ���Dj4��1
G�Aį֟CZ��e����OyHY��%;�%�Mѭ8� l;�}R�&�?A��N�F�'��O�zر�
*��-:A��(��R�i$�����D{��{�y
!��q0��w
��:���	��M��i��/O���X����m',"���/*al��eA�t���wyʟ����Oh��q�h�Rl�.C$~����D/��E�q�����?���"�3��в�¨� oؗ1R\I�A���M~֕�b,H�>�b��'�"}�'t8g*��~���֡	8H���@g�O����������S�>�^ �w��N���Cn	���'��N؞��]h�b$�'�R�XO�����<�	�]��]�	�?y�	Ǧ���E&*I�E�V�Ly�$��C��T��dX���N   �ID�'��-�d&M<	�̴�u癮Em���{�,u�����O��oY�D�'ٛ�%݌O��8*� �]&i8�Q��~�Mљ6`�6�O�$�O��O�	}�JY�$+��L,!�*��i�J���%cڜ����p>y�a v۬�]5���E���Xi:١aP*��u���ևIP�(ư���E|���~��R� En.��AOD�s�ֈ�Q/�O���轢��[y��'��'��ia-B-:!��c,��!@��)�{"�'� H���x�z��#nҰ(q�m�!	��q%��`ش�*)O)Z��A?� ���RmZ�~JZ1�Q��=J������	g�i>��I�:�������#c�Ηh�p�$�M:+qj�ӶH8lO�u0�c�o�ԕ���(���]-E��qAQ*]�lRe��ɳ.(,�D�O6˛*U��.Up<�rG��y���ĩ<�����S'X9�Q�S6J�h�x�oZ�w��C���v ��A��l�A�t��6L>�7�lӐ}lZnyr�Ԗ�6��O�c?��CC�dx���>T�q+�M����I쟴���5�	쟰%>�x'(^�)Ŝ���a�,nu�epT�:���Vi\�`�:J�j����)VHu�yՆ�<d�)������O$��7�'��5�I�~�&F�������.�@��e�X5n=�O���<QB��5d�z���X�|�浓�'x?q��I��M��i��4b�����ƛ�jg�}`Rə�u�MS� �;b�v�'|�)����?Y��M�㝿w�p��%Z�y�0�Se-I6ykE�>�*���>�O��)@�J%j���l�Q���iC
��8$(������D�Yv�i>�#}�'�X�i6⋿x�|E�B$�$?����DO�Ov���Ԧ���9��>��BJ��a����ү[�!��i��ub�	m�'�j̋u�Fl�8p���U��\я{�N`��Ym�M���rڴ'��b�ǒ��h8�E�Ȝd?,���+	��ĳi���'tr�|�O�fI[)A�8S��Ԅ)��-��Pv���7*�j��P#c 	45@�G�1A�����k`ӈ��E�N�N�J�u�'�^����*_PS��S�^h����T�
�����O�lZ퟼�'��Z��n��
����PJ�.I0��ќZ��B�ɲ �ޝQ��J�<$R��T�T�ls�,K���d���'B�'��;J�`�� @�?�   �  S  �  f  j)  v4  d?  �J  V  �a  �k  t  {  >�  <�  �  ߙ  -�  p�  ��  ��  M�  ��   �  ^�  ��  *�  ��  �  H�  ��  P�     L � t � ' �/ ~5  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z�����W��K�L12$���SO�\1Yd�	�O�!�WR�H�Ī�.b�&hb1[��Q�|���T>�%		i�JI����z�`��6#1D��Sea�d]`b%�\th35D������?!�-Q�ė
?<��F.D�@3A�	5�Fy�B@WD&�H�!D�,s���CB>�rR�>dwA�*D�$0R�Ō*���B��30�)�-&D� c3�jFM �jp����('�ب�^��*�\�Xi��tU<Z "OlA�g`�$`&�@��I�kHH\C#�'ў�
Q�� P���]>�h���$D�\��.�h���p h�X�\�L-D������~`&A��K 1.V���5D�x�`ך_s��:��Yd8�4?ю��S7\�^5 A�ݯ�R=8�'��B�IP�&D���� �DU� �#$��B�I*1	@��G���J$E��LOO�JC�ɨp�\Dhfe�?`��鱺@�e��=O��i��b�x�Y�)[�ks$�ȓk��b#͔)rNQ��K�j>-����@�w�B�[*�� G<@�-�����DNA�R}�U�$���g\�܇��i��T}���.Ƞ��ĩ�C�(��C�	\?ы��?vԠ�F��K�#=���T?t���N�\Ry��:D��ۢ�b0t1��,�'b�tg8D����d�M{��CK,h�����5D�g�7Zr�#�o�!}�%3�B4D�pn\t���V͞؎i�sG0D��ڀK��/��r"�0�r%)��.D���u#�l<���`��MfNݲ�M-D�J���p���s�mX�1F�K7,D�PsC�Rj�����RLmXB%D�d�5mc�D��aiT�u:8}��#D�Da�H/6)bY�dݹV(Yxu�-D��Ԇۜ��e+���
Z�H�c+D��c[1N��A���5���R�j-D�xJ��S�u����@�b�``���,��h�4`Gf����B�f��C�Y�h �ȓ&4e�R�:�t�Bt���4!�ȓiW��
G��#�>L�s��)�z��ȓ3��Ց�B�	N)��ܞ.�4���o\\x��63X�p!Q��2����r��)9V	�4!(�E��
yI0��ȓN#�S ���(HG�ϭs�b�ȓM�@�y��/^��6"L�Q�ȓT��"��԰�h���֡�X��gX����H��O \�j��%g��ȓ.��0r��ݍ4�8�Q�<o]
@��I�L�Ӄ	"&^B���ǻ)�r���<�@,h"�L�\.t�%��6���+݆=s3��W���!DK҅��݄ȓ�z(��k���V��EU�j0���ȓ�R�Z��L�^��+��Q�k2(�g��~b��Y2���Mۉ\�����[��Ov�'	|�c)�*P�ӋA�1��Tr��,|]
g"O� t��v��,l��A�i�#�A�R_����)ҧ �`gc��Qq��a�.Jž�ȓT��1ٶKW Ĥ��@Ж3[^�%��z �'���W��-�:P�gK�.�p�'��Vhe����ȝ����9�bB�ɚC'B$XEi�3Q���R�( ����RO�tJ��BЅV�h�k�$G�n���BG(�<J��C;c��Ӳb[7L��09s*LO7/�I�QT�b�-��,r^ѳ'ɍ3?�*B�ɕ{�z�12LD�|��x9r�e�RC�I�f7�a��`� }�D�����B�I�5cZ����P9��S"S�84�"<�:��A�����Hy>���M�9#.�@�ȓC|��+t�/)<e@C��7hL�ȓ~��)��X9{���R��;'�<ф�J��,E�F)�prc��r���ȓ&e��[���88�£�8Mu�q�ȓ]o���1(�v�z���0rp���S��,�?W�Rqj��0)���ȓv�
�p��<@��x�t�������{Q����nU{��@�FF�����J���7 J%M��1)P ԂC�Fź]�� �5ݺ vNQ�a]�C�	(,�x�H �+��PC0!�)O�xC�I�$ޔreM�]J�s�OO�%�C�I��
��
�;.b��Q�����@B�	�Sh�H U��2d��vޟwu�C�ɐE������ ,B�2aA��j2xC䉏*hTŁw���x�ʴ�Z�}NC�	=<a��j�#9ZB [,W*�<C�I/odٚ&KиO��32j�>C��妰pb�S<(�6���'���e��&Pb���+ƾi�0ES���|m���Di6ʄD44$�[�oI0�^���>͌�*R���+�,�$%`��&v��Y�G�D���\�kڦĆȓ?8��(p�-^`<E�.��d��,��2B�ܻA������=��ȓq�*M30a B��r�
Ѭ��ȓ4ᐥ�$�G� ��u�s�x�\͇� xp� !�\��Ӆ�f����\6����?O����L��$�\�����I?e����$BXQc"O0�t��~�����L1}0��{�"Of�����x_y�3mυn(D���"O��ue� .��AQĂGT�c�"O�к%'��_�� (��N�;�>-)�"OT%���N=$��0f1=�Zغf"O�3�ɒ�}��%E��_��5"O ��g̓��V}X��ܖu|�1�v"O��h3�Ɨ$b(+����'U�)�"O���p��E�P0���s6�hA "O���1���!?@P��ͽ[���"OH�	c�$z���q��W�hXX� �"O�,�!FL��`@� ˭0@��"O���H��"�:�po��>:�""O&�h���Uc@��w/�uS�"O�9���N0�@V�r p�0�"O�K�b�g���9WE����	�"O��@��˜txs��u���:�"O*���e�j&ਣq�Ʌ:�xa�"O�X#`gE� & H�%�S���:�'�u�aL�ބ	������6D��2�gX�Fl�!�fG�5N��e)3D�� xk��+�:��Ç�'���d"Of%k�߃3s�l��On���"O�0;r��(A0E#�Í�5VΜ��"O��炍S��(� ��Er��J�"O�첗������*ݜA�Z-���'3��'���'b�'2�'�"�'=Ҹ���O�:�
9��pxF51��'V��'���'I2�'���'B�'X�)�w˗�c��] �Λ�c5��0B�'���'��'	��'���'}B�'���[���,8xT�,ݎjڌ�4�'R�'�B�'qb�'.r�':��'}��[ 
жO>^ԋ�6	��P#�'�2�'�B�'5R�'��'���'�0T��ˎ�uW��a�h]�0�4=���'���'���'b�',��'�"�'��\���l��Fj��JM��':2�'��'��'��'���'�]C@��'k�����^;P�����'9�'���'T��'H�'���'QlpZ�D���'���l1��'"�'�r�'+��'��'�b�'x�U�As}�IE���Z����'j�'ob�'��'k"�'�2�'d�ū� K;6\d�C�[�aNİ�e�'4��'���'!�' "�'D��':43׮�Q���jҋ�"dR����'�2�'�r�'jr�'���'Xr�'�8�[W�+&WV}c��C�H0��'���'-�'{��'���b�J���O4�I�;'� )��ܒW�L	geCy�'J�)�3?��i��M#Q$߼P�\�8T��4p%��۝'D�I	�M�R��>���`�䉈c���Lt�q�����
��?I�&��M��O��ӓ��I?�f�ޡ]�Ѐ!��_)�b�f/�ԟ�'��>ũ!��7��;ƯU+
n��s����D�<I����O��6=�QcT��� �z����:Lbpͺ�"�O��e��ק�OG|��i��$�8eђ��9@8�YWEL /��q���uUƢ=�'�?If%Y�0��&�;K��`Պ��<�-O�O��~��g��!GҢʂ��@�	�mS�2c�>���?��'��ɷi��(��K���#�k��9���?�ă>s$��|���O&����Z|����De�J�#W�'`�U�-O�˓�?E��'Ij����;�
}�)Ij~�9��'
����$��9�?�;Tb2h��� JM�`k�Cݺ=�����?���?�pe��MK�O��S$� -@.� �H��\�h5N�F@�
?# �OD�S�g̓Ħ]� �9q����������'C�ꓚ���O��?F� �nn�!B�����9Õ����OL��9���M�;v�|U�ȉb+R(N�H�l��@��U���D[�M�&�O@Y*J>)O�r�`� SF쁶���ļ�;���O��$�Oz���O�ɯ<a X�\���t��Qjt�ܻ<f�X���D������/�M+��>����?���;q(�!1c:�ȣ��]$J�j��W��M��Ot�X�ʀ��(���4(H����ϑ���"�l��-�$8�O��ꅍ݈P̶)S!aR�+��Ai�<���Ss�)ڷ�i��'7��3��DD�X�,0�P!�!VM�	ԟ �i>ug������uGʜ�4&,`��ေt0X�A�����[�'<'�ؗ'���'���'�9S�+?0�.p�&V��r	���'�"[�D;�O ���O�D�|�!�!+�x��C:��Q�`x~"�>Q��?aH>�O���c���
��<����621|�:�-�.&� �B�i$���|*u���t%�H�̌7c��%�CȒ��3&�ןD�I۟,�	�b>�'#�7���I?�e�Ч�wL ��>.��D�O��d�����?Y0Q�����iC��yu��+T�PX����6˞���ݟtj�cæ��'w^M)*�?Ť�܌YÁ�
x�^������t1O ��?���?����?����I�Jtԝ����=��Uq੍�/�y�'��'a���'M�6=��)�YY��1�
�iu�Iic��O^�:���ʍ:�6�p�@�Ư��0�p�v&T�^$pUh��m���c��mc�E��ty�O_�Q�z�{�(ȣXw��ht`;_7��'���'Y�	���d�O���g>�!��X&c�2���xU3��+�	)����O���)�DȫP�qz��0�Z�{�[�D��ɣN��ٰ�����|R����ɻ��u��dC^�Q���~#� ����	֟���r�O�Ҏ�z�J�����8ت]}�""�>����?iV�i(�O󎔽{��)1̂�E�0�$�7���O����Ov����w��;��� vG�?���`��2��pH��� �h�	Sy"�'&��'QB�'��`��B�vK�$�wK�t4 �S��	�OV��On��(�)�O���&�0Ӏ��ܵ4�Y����k}�'��|���J߿<H������'="*�����d,`^P�"���OZʓ^��a`�M� /g�
ņ�:I~���?����?���|r,OhI�'�2BD�3H�R�р�\������!£f���p �O.���O�-�	���1\ǜ	A�*G�G�h���yӔ�y�I@wK�?�$?��=� ����%$t�zP�U	L�e2O��d�O����Op���O��?��A��B�vi��!�~��}hB�ڟ|������O��>�M�M>���]�8H܁���,=�9��<�䓜?��|z0��$�M��O.({U�ŷ,À�J4!�w*��� �E��rx��'��';�I���ڟ���62Ƹ#��]�)54�B`jC�B-�}�I��4�'\v��?A��?9+�Np�rϽu��2�P�2��iR;O���k}B�'g�|ʟ�8�B��j@L�2�	�HD�S��ԦyZQ"k�`���T��K?qH>9�$�PqpD��U� ��p�B��?���?����?�|b,O��m��X����+g&aH0��d�F�	���	�M;�B!�>1�s��	���{���0G�-8LP���?���M#�O���ea���P���34�*A(A�8-�e�`�,�'8��'���'y��'r哶2=n��ˡ=L���	}vҭ۪O�d�OR�D:�)�O�oz�c�!�:n$S�]�j���S�П���r�)�,�n�<I�	Q�7�0��f�6�����J�<i3MHih�$^.����d�Od�d'(�Za��k�K�hPacd�/j ����O����O�˓C&��ʟ|��ݟ@��+ L��XF��@���U�8`�	����B��
���ȄX.|���è	uC��\�-��@�&�Mp��4āA?q�,�ʐ&ƜX��`��Y�S�8�K��?	���?���h����� ,�h��R7R��
���eB�Ą@}b�'&BBb�N��]G�>u�4�-
]����3J���I�����̟�hbA�Ԧ��'3p���R�?��4&δ�;"&�8&\���H�6b�']�i>���͟��	ڟ(�	�xW>����;w:B ql�Ґ�'ߠ듡?9��?iO~*�������I#S44h%�߫j��-9�[���I��t'�b>�&��9 ������䂀+�)Ov�m�`~��� �>9�������;V�\*�f��G�p��L�-%TN���Op���Ob�4��ʓ7"�	���ϨLh�Ɉ�@��1�V�h�8�ٴ��'�N��?a��?��:B����Մ��(��)C�|�4��D�!�����'f疓���N_�����X� �>%�B	�"p�d�O����O��$�O���3�#sB�\0!AաQǊ�2�+�[O�<�	ğ,��%��4�"���M&�d�TB��x��(0dQ�u��0:ECFt�I�0�i>iac˦��'�,EP�IN�~+�@�����9[�i ��¼����&Y)�'��i>��	���I?�( ۓ#N\ЈeX֮Št�	��4�'.v��?Y��?�(��kj۞3�.`bn�0u��\r����H�O��$�O��O�
��E�LL�36~�*�Q�A�zu��\��Z�ls~�O�\����%.5��*�?X@`��6 S^j6����?9���?��Ş��D�Ʀ�3t���/@���L���؁�g����ܟl�ٴ��'{F��?i�&�Rʀ5�WA�|�>��˔�?i��ed�޴����2w��Z������Y�0���(k&x=�5�ˈ�y�_���I|�I�\�I۟�O!����K	�G�"��C.M��y��>���?�����<A��y�o�9j�Y0&	# ~���5&P�RX����D���6�j�pàS(Q�앛c��
�r�h�*s���ʞ�8�)�M��{yr�'��Y�	t���I�<W	 }�p� R�'���'^�	����O���O����e����y� �%Zp���*�I���d�O��D=�d�l$�����D�N�B�鞿Q=��%���".^7��-'?I�R�'��	���X�\��1ᇳ>�ƱKq��N����ڟ���ퟜ�	b�O���G?U+TA ���f��=�煘�-&2��>����?Y��i�O�#Kf�L�/.?�h��QT��Or��O����~�*�Ӻ��7��d&�\�r�+qƘ'[����-�B@�O�˓�?y���?���?��R�P�����e׺5�3�[� ��/O���'��'���I�=b���P,�+n��b�G_�4��'	��'<ɧ�Op���,^2'��3��#dQ� ��q�֋�<!���J���Iu�eyr*W?:��2��'"m��a��'PR�'d�O��	���d�O0���P�0��P%��	9L�O�5m�h��r\����ܕ'>��/v �1�/:�)5�!L��р��i��� F�0� ��Od,$?���#:�����P�-:��cb�I͟,�I̟(�Iן���H��dNX0k�gKQV���a"aurpc��?Q��$�i>����M3I>!�n��~����a�
g��I�7���?I��|����.�M��OJ��f��"��"��ՋcJp�S�Z�r�.9�'��'���韬�	�� �I�I�Ķ6�jh�ɣ��[:}s
`����ԗ'؈��?���?y/�
�{� G	b8QBa,>)�hӕ��*�O����O`�O�ӛ��T��ˈ�|,�� �'!���0iO�|R���W�<?ͧ3����C9��t> �WĜ:8\���  �	�����?���?�S�'��d�Ҧ�	7V�eN��Q�-wܒ���)c�D��ɟh�ߴ��'����?���P�j���J�	o�m+����?���q�`i��4����*����mk+O� l!�s��!`1^�����g^��9O"��?���?Y���?������<���P!�}���`��(�xh�'<�I��0$?i�I��Mϻm8Z�Z�o�m��	A��Y�b3�����?�N>�|ʷ��M��'�X�ZQ@�5�(��DȄf��q2�'��Zc˂��dhƙ|"[�t�I��l�T" 	���ڂ4��Q+f���h�I����y���>����?��ф�qį�V��R�(�<�@A����>q���?J>Auj^2�6�9!���7�P�R�K~bBZI@�I����OB��	n��+P0C' bfͺ:rN�9�-̉j�2�':b�'���S���c��i���6Dͷv" ��6a������O����O��mZ]�Ӽ�iә��"���-��XFh��<���?��8:����4��D�-:֘z���u��B4uT���5��M{dƐ5����4�����O����OR��n���f �2.��>	���D2����I��&?�	�q���b҈�'{���*�a�.H����O|���Ov�O1�Ԥ���a$��c�Ӝ]�J��2J��*%�Hv���
�`ԼUP2�Zr�}y��?��`�y`�;d�C4���'q��'��O�I����O�,z�lV����!p� ,����M����Ħi�?�P�����杚^��1�4e�%7�T�9��P�E�N=�B�Zަ��'s�;���?eY�����w"�b�@�3��Qi5!�9����'g�'\b�'K��'��V���'�"�xY�O��-���p�	ҟ9�OV˓1O���|�0 �ưX6(� � �B��Ø'+BU����U���'��������^
K�D|���M=����'���$���'!��'��'s2,z���\e�s�T�(�I�'�BS� ­OZ���Oj�D�|B6�Ј;��j��$+qp��V�X~�,�>���?�H>�O`����O�ډ�cX�B�XQ"&έpsl�ˇ�*��4����Q��O�I��˻���p�7�rH�I�O��D�O����O1��ʓX���@�P0��#J�4}4�A����yB�'3eq� ��ѬOr���'�lUJ�\]���S�+#(���OT��c�m�,�Ӻ��ޓ��S�<Y�O:˞}cрˑhb����%O�<�+O����Ot��O����O�˧k�� ��
>�� 	pN	��p0PU���I��8�IM����������`GL53ۈ�ׁ�0_�����?1����S��T��¦�����YH��W*�"W.<%�FEC7�y��V�z��!������4���$�x���ՈM1@�`ʄ�
6w�h��OR�$�O"ʓd��IKy��'-0�]8߸��ѯ�W4n���|b�'%L��?����H�ʥ� �B@��h�j�� �'��\A���NS4 ����D�@�(��'��A8u�P-:Y��Q�_�a�I�����͟0��p�O��#G�$T�y���>�ԅi#d؛t3b&�>9��?���ie�O�E3;�6�����.��hE�9_��d�O����O:ݓ��b�v�3�DifN��� ��+�t�X"�4	� A��\2�䓞�4�`���O:���O���j����j� �m��F��˓K~�	Ɵ,��ҟ�&?%��3֢��� G>��g��\e���OX��O`�O1�U��� Q`n��ED?8��18�M�/Ȳ7m2?�� �,���M�IWyҬЮ*�:�:���C=<�(��΢n�r�'8��'M�O��I����O�����"(��@��=QGt8"��O�in�@��u��	�h�	П��KN�C~�Щ@��y�V,�f�ٷ1ъ�mZc~��g�n��]ܧ�����3^dd5����������<����?���?��?y��d&��>���&Y�s�=��Ob"�'a2�>�'�?Q��iB�'&~��q�"+mrh� h �]y�Ĳ�y�'��Iq�BLmy~r�Gm�*�a7g��+�keh��#&^�dq�|rV���������ʟ��Р�q�:A��.T5E\wc�Ο��Ipyb��>���?�����F�&~�L:��L?x� <sD@�|O����D�Oj��+��?iZ 
�q��xR�[8���g�����A)U�'O�����$������|����F�8YǍ�
i�����I\s�'���'����[�l�ܴ��*��a�0���n3�f]�<���?	&�i��'m�>����d�q��vYj1�԰����?A��ߢ�M��O�N ��x�I���$V��T��==a�Z��4)��'@�����	��d�	Ο��	\�T���}sl��Ւm.Θ�2��-Db�����O䒟X�d����/#�g�ƞJ�I����nh�x��ȟ�%�b>M��A��ΓrDX4IG�^�*�X}�2F��X͓udX�"2h�O�h�H>	*O ���O������3�RYP��%�.���O,���OL�d�<9�Z����̟T��/#*�K!��*$��A��iڝ|���?��^����ʟH$�x�G�O�Y'��4.[�Cw,a��OTdʕ-�V��E��"�)F��?����O:����m�*�j.]�^�6 c/�O��$�ON���O��}��^� �cZ�/�����"R�����	ȟ��	�M���w����NV�-��'ڳ:0BpC�'�b�'p���j�v��ĉ�����4�>� \��D�K���vh�Yn4�A!��<ͧ�?)��?a���?�'��R��{�Ġy�(p����ċx}��'���'l�O�d��)}��Kƛ; ��c��0`D��?����Ê;p�XR̕��ܱ���-3A*̨f�\���?w��(�`�'7p'�,�'�p��΂�)�.m�#P�%:�� u�'�b�'Z���O��	�����O�5�͇�=�xX ��5#��|��O*�mZN��n�	۟�����8����ME��b�L�hLfEȠ�A�t��nZd~!	��lD���w�Ĥ)�	j�)�Cգ#	�(��'m��'t2�'�r�'��>)�➓�N�G+	�f?�qj�<Q��<�i>�����M�K>i�넔{u���bʪ���GK���䓲?���|b�W�M��O뮏�sԤ��/Ҿ��Dz��ʲ7Dވ�g��O6�I>�/Ob���O��D�O.1�P�XT�:U�"&*,�,5�v��O����<95S���'uBY>� ��F��rx�GG�/���g-:?�5Q������$��'�Ҍɣ@W�#�Px��H.O��<��(�����KDK~�O!hI�	���'��ݣb�?a��A�p^8N&|�v�'xR�'����OD�� �M[`S>]���bꎉӖ<���<����?q �i��O\L�'+�m�3h�+��ZnЬ�����'��g�i*�I�J�cq�I��GZ�(��~�F��ƅ��K��<���?)��?Q���?,���� �
�~?�!�g�4Fʈ9�O�V}�'y��'��OxRdn���!�4��!
� o�q�(֯T���D;�)��06Lao��<q��l�ܓaA�<E��G��<���=��Q8����d�Ot���&��p�LVK��ェ�\����O�D�O��r�	����	؟$!ҫte�BT��c��9�
@-}E�OE�'!R�'��'QX��0%�6T`�Lإ�S�!$��K�O�4��_�Xe�py��,�?)��O�X�������ܼq�,��en�O��d�OF���O|�}���'Cr�)��Z�(zTL,U����Z���⟀���M�M>Y�Ӽ��K�aw$(���!Q��Y���<��?���r2�1Pݴ����R������Aa�K'W��0c��:S�ȗ���䓺��O �d�O����O<��A����WK�� XS�/Ԓe��ʓ)0���`�����%?e�I5s���xF�72f���/];~PDջ�O<���OʓO1�ִ����V̫�@!�`y(`M˱P��7�+?��a��(�D��J�IUyr����} ��u_bD	�	�+xJ��'�"�'��O��ɐ����O�M��ݼjC�!�$��CT�L
���O��oZr��p��	�X�I�ɰ�Ӣ{����B��cK�l��	S�p|�-l�a~��*Lc0<�E�'���E�fN^94� >
EP�0b�<a���?9���?����?���$d�{�oЅ�^��ah�e[d}*O&�d n}�O.�cr��O�=aU���h@�Y\\��!�+̮z��'������<e�6�0?9�S!*1f��a-͇!��)Q�GR�M�<M���O�|J>�*O�I�O��d�O���M��@�ҟ5;�P	�O$�Ļ<a�S�X����|����cƇ6��"�ӱ>�0@�����Dc}B�'��O�3���$M׌;�	B�]/e}�t1��؜v���Ry�Oxb��I�C�'� P󂓼U���
ˉ\p$I�'y��'�b�O��	
�M��l� A�"�� B^@�Vurs�E�<	��?Y��ie�Om�'SB�QGyD���F�7M@�4c1�' 8y��ip�	Q\��Y��I?Z��m�5Q�_
x
%��G�<Q���?����?����?�-�h�� ��.��0r/ʅq}�(�c�Pb}��'Pr�'���y�es����A�b}ӄ�P�Qh:5�P�$�O�O1�v}�Kl��扁qs���t�0 �m����)W�物J-~s�'�θ&��'���1���	�Hϵ��ta`JPY������w}�U�(�ɯ8���C`�_�lh¯̑o^���?9�\������ $����%�5Qo�h0l�`6	T5?9� ӌG���˖��O����?�Ǥ<fQ@��-A2K�4�BSeĔ�?����?Q��?y��)�On�["�*|���Tk��iWd�OY�'���'�7�0�i�q��e� z7,����!��y)gh����ڟ��I\��<n~~�j�;pQ����������� 0B0[��:��u�a�|�[����������	���"$�c9v�zGOV�;�X��c�y(�>A��?!�����<�dőE;<��b��B�B���#�YG�I���?�|:Sl[CҰ3#�- ]�D�G�<���2����$&�Z�c��4ΒO\ʓ&v��p��_�,���+��xJ���?A��?1��|B.O�'I�e����Ӱ#� ;P�d]�X"	�b��J�O"�$�<�`��FͺtZ%�O�^`�!�o	�/�����4���ľ>( ���',�F��8��τ4����@\�Z5����*P���O����O����Od�$"�S�{�l�h"�˶{H�Q�ݕ���ɟ\����$�<�g�iW�':��1���A�Aq�.�5�\՚�|��'-�O��9P�i}�	� =�� R8�5����(C��&����#�? ���<�'�?a��?T�@�3��<p�D4g7P}��C,�?����@}B�'�R�'��ӍW���J�f�fy���U�]�v�|��I��\�?�O�h|��BOgN81YA�윳��F�|v��Ē
��i>m��'N*&�T{@��?r���$A�;��Hc�P��|�	�����b>��'�b6�K&�EB �?LA��e�Lm�<Q�i��OTA�'�r�Y=x�x�v��4p�f�y�&��C��'�<A�i����&��M{`�Or�&��DBΔc�
삢��'��<�,O��$�O��d�O.�d�O6�'>w:V�E�&�� �V�lP"�IR}r�'=B�'~��y�Ga��nܭ~��aH�*l�*Ex��Y*TqF��OF�O1��UX�r��ɏ\^�(*���e[L�"v��an��	�'��I��'}0-$�Е'
�'�P��$�{�R�"5���{�>T���'}r�'��X�0	�O>��O"�$A��~<ӶB��6�䭔O��z�O~�D�O&�O ��w��YZ<��(՘o8�����x���<O��pq�'3�ӿO�'S��JQđf�ĨH#oDh�D������ٟ�	�DG�$�'�*0Ҳ U<��3`�6&z����'=.��?���S���4���(Go�)OodB���b�DR�1OF�D�O(�䈥p`6� ?�D��4�����M�D�8��Y�pl�К@ �4J�8�%�ؖ'j2�'@��'�R�'�@���B�T�Y:��)�l��_�T�O���O��=�9OI �,1��ʦ��m���@}"�'�2�|���MM1V�3�#�)�-����a�:4s�i�dʓ���!���$�@�'���PK���X�%�Q�<pRB�'���'7����Z�p�O&�DZ���I�`�L$�*����o4�D���?']�T���X��'e�4��TH�0�
���5l��Y�CԦU�'԰�B��	�?-�}Z��S��Ab�H�Dt
��OC�IpΓ�?���?���?)����OnDAzTd:?����
�	up�K�V�������4�����٦�$����1~L���[�x��cq`Jj�I����i>��W�AӦ��'�j4;��P-�łD�cQT4@7��8!�l�I�Y-�'��i>��i�MS��`ʜq3 �VcF�b��5Im�����?�/OFM�'N��'^RY>�j"�I�5lpzpꗬz�,Q �e�H�ɤ��d�O�����K$�Q�!(n�ha䆋d�p�!W�D��@��C���'��4+��!��|�JQ��y�GM�W�*�K���e���'t��'E��4X�hbٴtf>�s6!A�K�vEZ1/�6�����?���v���|}��'*���#
�v�p�%K�v��M���'8�A@>>�摟֝�r��Ӝv�割>�D���o�QC��R~
�	@yR�'���'��'��[>�hR	i�|���5|y	gA���$�O��D�Op���������1o�<��� �)2H�u�2�v��ٟ�&�b>ᑵ��Ӧ�ϓ4��(  �	?�"�Y)z� �  ڜx��O��䓄�4����]�Xr$��%��-�zy(p��1eמ��O����O,˓@��I�T���|)t�-���kV��-iC�W��5|��ş<�IX����(�L"� ��O4RSF�E
\A��I�Y��@�|:���O�@���Jq�j	R��1�R�I�.���2�L�O4���O<���Or�}z�� ��c�N�wd��6��&&�j��xg�Ipy&{����:`br�� K_'	�v��v����I���	˟�yO��)�'.��p��?��a�ܤJ��EO�R�JU[��I�l7�'��i>��I�x��ğ�I�>���$�~�i���(���'e���?!���?�J~Γi�\�#���v���lު!$=��^�4���%�b>�O߁$S�p�׾<�,y)�e�I��>?�R&���<�d
=����	!|�b��sm^�*yv�i�ҝy���OH�d�O��4���!]�	ҟ�fl�b�����>db1xD,@Ο<�޴��'/���?a-O�R����ar�嗿	��&�Ϗx7M!?q ���p���iD>����V���ٳ�ED[�t�m�!�y2�'�r�'��'r�IL�v�!�V�; ^Q�E�����Ot��j}"V�X��4��B�l�Bg��>.1�<�u�ŝuF��	L>����?�'�� ��4���P(3�`�DB��3ڬ�Hu�^���D'B&�?i��:��<�'�?���?	G��;&�P�3��)��[&V��?Y���D�W}��'���'��1�D�r��,Zq<�C�	[	���I��Iٟ���b�)jt��Z���aJ��`",�:��RF��7MSk�V���ӮrC�@�6��-*�Q�Q���L��\�e)��|�ȕa��6�1���*G�ʹ`�M�J5�X�}q4���+� �̑	d�K����E�?l�b�*ƭ��b��ׂS)t�����-.�K�]H�Ξ
J��Y*r�_�0��=��)�������R�����!�*�[ ��"O�H�����; $a�+��3L`�S���f�06��9:���4G��L*ŬE�k����3I,s5lې�ƩH�Tڷ�X�4����B4 Ű$s	ιg�fm�p@]���S샋T����
&C�:�@B��*i?���>,O��D(�$�O����3)�RM�V���D��C��Jx�*�O���v7O����O��$5�ɤ?� 4�2�DH�y�1��Oh��H��iCR�'��|B�'�8`Zc/L1a�"_fPh����~H�X�-k�����4�	���'9����4a��W�~��"�(�3n���f���M������?��cNT�a�{��J� �$��� 6p�8��M���?��+��<A�����OB��O9��F��iSk�!����Ң�G�����ɔk�r��?�O���N�-Ee���&�X� ��4f�<T͓�?����?A���?�����ٸ9M�����P�|stI�%4���n���	��nm�?�O%�0*�4cHʂ"ۄ:�$<@#.��l�ϟL�ش�?����?���m�	Dy�CҿR<���	�g��c��ņ�F6�����D�OzH�'��ē+T�^��^��68��W
6��O���O��A}�W�(�	}?!vN
�aP�5�B!ά3�"����FX�x������V�x�Γ�?����?��dH ��h8� "�h�&�M�6�'G�>�/O���5���<�{��X|�T]i2 ��M\0��R��7J�ҟ�u��|�	؟|��f��H!p�v�у-[OyR���_!���ly��'�'k��'@�����2
 ��ӷ�C1q���kCh4�y�-A��y2�'��'!�Ol���E������j���V(E�:��7m�<	��䓗?��7-r���'3H5�"�L�E��Z���lk�L�	���	��'���Op��My�`$�,��^�ؤ������	D�	ß��	���=���[��(W�_/%��������Iٟ�L{������	�O����Okǧ��%���:4h8�%�A�cF�'t�	�L��L�s���!�� ��
��zrT�S�	~6��_���Oh�oZ˟��I���	7����3jq��qk�'6�Z�H",,�V]���I���aI|z+�NM��iμ��`n�`s2%�!m�k�D}��'��R����KyʟHH0fY(��Z�FQ<iG�` �W}��%�O󩎃��ɾ�𥱢�N��=��]���"ٴ�?����?�����?a�OH�����S��Y�w� &1��qk�_[�'�"��z����?�Ӻ{����1�r�R��:D3"�[�IĦ1�I��|�'� �'��'�	�GǛ;��A�cһ>"t�Ƨ%��ҹ5��$�����S_?��C@�.!�h�ӗ6Hz�!�
��'�2�'�Od�Ģ���2	�*`h�4;��ľ o<E�Fnt��|���.��	�X�i>��'���r�P�
�F��Z�XM��ݴ�?����'W2^�P	�&dӐ�3�`�/k�Nq�)I��n@+����<����?y��M��O�8�'�?!� �b�Ȭkc	0�%+��Zm�V�'��'��i>9�	B�	^��^Ţ��Z�T���Xw"GvW���'b�ʇn��E���'����56�M�[B��P��(=>�m��ē�?�/O� �u�i�U3Qb� �2!h��(�n�8�FxӶ�[�;O ��
������$�	����O��`F@T�ZY��*�d�i��`�7�i�����I���'��� �EÛ��iOt�2�.�!T0��`�n���D�O����OF���O�S�Tc��X��lޑ"�y1$�&Q�0�p�Fx�OR�ʛ'��(�A$P@#�
B�6d�!Be�"tn7��OZ���O(��m�)��'��IKhH�/'��X��5t��,�ݴ�?!K>)����Γ�?I��?���_����A�d�0��t�s�7S����'���=�?-�'��� Q2�!v�-vg̫o��'�R'�y��'cB�'��'')�I�b.A�~)��YA'���2�n��ē�?���������dj7��?2ZuA5��@.�� ��i�b���y"�'=R�'H�O���S��\��$�+6~�� �A�^�듧?�������4���Ē6���"�طx_��J�;FWN��0O��d�O��$o���I�O���C%��T����hY�9���æ��I[yR�'l�'-Dq8�O�i����C��Ѕ�w	T!$!��4�?9�� �|͓�?1rY?]�	ğD��/JE�P2�.B̙Y��T�x����O*���O8��&N����O�ʓ������e���/ �>L�c��	�M+dM��<9�x��'���'�Bm�>��]:��qD�%T��"� �d��o��l��}��IZ�Ij����M���L�'7؍ �ж[�hĢ֊Z��y���M���?���?Y7R�Д'_r1�t@�.]�0��!��2�R�}��	�<O0���<!(�ƹ�v<�b�D��J��Xs�ɴZ?���E�¥0$o�ԟ��џ���=��ĩ<���~�̖b�����=r.�M�u���Mk���6��$� ���O����O���h?2H<��TwG1C֏����ߟ���O(ʓ�?Y+O*��ƐDZ�-�6����獤(����_��D�}�����H�	ȟ<�	�?�i݉��gXz�"��aCͿ:�����{��'>�	P�'?b�'	�J��V"�JS"�5T��H����o����'����'���'<2��$�>y���)���o��!�,|�4��?�/O6��O:�d�����1Jڢ\�fI�Ch���ٻcE��X��'W�'7��f�m�O�n��?�1��Т�H�쮁��c����l�ʟĖ'���'+�/�)ߘ�M+`Hϱz�ʗ^#�=��/U�H�7��O����m�D�O$�O���'���8� V��$LbG�TSiM���Qf\���ʟ��	���	sy��'���L�/p��0H#2�ظ脖ś���y��'�7-�O���Oz�`}Zw�SD�Nd}{V�C�kV^���4�?���~��������u(��$U�g��R��Xc:$�ed�$�M#��B�6�'A2�'$r,�>I*O�<�(�!����.V*�!�B��Ѧ�X�%p��	yy"Q>�92�z>����C��lanӚa�l����e�V�ٴ�?��?��&!��Zy2�'_�d�3t���Ȅ1g���Ӷ�+_���y���yr����t�'���'��*A�fz*�A��Ǘ�>u0��n�"�D�O&��'v��ޟ �'wZc��l ��a�0���	p�D�@�O,�&2O�}��%�OD��Ov������B �ν1�sW�do��d�i�f����O�˓�?I��?�/��}�~qdT�&t��kdfE2"�Γ�����?���?yO~3�����-��EDN�a�#�)h*��V�x��'C�'���'�Zՠ��'߾���2D�5p���e:��*`L��y�'���'8*��4�O9���=y����Ǐ�-rݸr���pP�7m�OړO��D�O�`�2OH�'<���_��v�y�!�Sֈ��4�?��LP�͓�?YV?e�	ş��1cLL{���2�܍��\�`��N<���?��b��?YN>A�Om�,�GM̫t�5�R�W���`۴zVt��?źiB�'���'X^�U�Ri�q�J�YQ�� �Q!Sr��m�X���
�x�Iu�)Bq��Ӧm{����	��0��Cx����z���WզI�Iޟ$������}��_�L��S�j���Ē{�B7m�'&Ph��#�$�|2g�R�<I��i&�͑��+5Q�I�AD؜#�as�i���'=r�'��Op���O
��O]昳�? �]բ�=o�7m+��ژI��D�	��O���O���aO�*6S�1��.N^Ԙ$�͝���I��$�K<���?�L>��*� j�D5|D����4�&��'�؈82�'`X��'r��'�~R�-&]Hu���2�̆Ҧ8J<	���?�H>��?����� Paǋ�\b�囕IT9P�Щ��j�B�ϓ�?a����OH��ST��Asr�S�9����S�P,M���?)��䓡?!�y���x�Z�X�b#�
6��A� Kk��¦�Ҽ�y��'���'T���h�OU��p��a��^�I��dx��,��6-�O>�OH��O����:O�'D=��(��^��3.�&���4�?Q�I�8xΓ�?9W_?M�	ʟL��{�m	`�S0����;v�<�!L<����?�g�H�<N>��O�X{��ÔIҡg�D�i�t���4pb�ϓ�?��i���'W��'Ϧ��0Y�˜<h�^%+���RE^)o����	�ut�e��j�k�����M��A��P唄�U�Ʀ���*�M���?1���?�x�O<F�0��7�ƕP̚�E#$�[���>�������#E�yr�'�����
=Z��&��(&���jk�����O����O�`�'=�	��,��r�:V�U>(
L�1����9m�ϟ��'{����'Ƭ�P�O��'��#�%ReԈ*��ŇJ��x�'	���6��O���_}Y�p��Oy��5ffS����@� .��������<�D0Og,�D�O��$�OH�9O�", ��(u�Fm�P%ߣ6{���>	/O���<���?i��2ۤ��w��m1Hْ�� �yۨ6���<)�lK��?Q���?�����)�T��'6�li�+,J��AM�eWNxm�SyB�'{��ӟ��I�D��Bk� ْt%LAR���9M,�#LT��I�0��ҟ�3O|z�Y?��It�9�Bl�<[�����CZ�ՙݴ�?�,O����O\��ٸSS�Į|n�Iʡ�A�0_�P������-g|6��Of�D�5o����OB��O2��'>�������xr�n�lAp�f�Q����?���?�C�J�<*��d�?�3ƒ$b�Ɛ��V�n����v�>�i�3O2��ܦI����I�����O��wJ��� �&%�E��&F
8���'���Ԫ�y��~�������y��΀�0��h�"��`���󲇊�?��?)���?y��?�*O��ER�H�'�]8y�IThZ�=R�\K�O<4p��i>鲣�e�p�ɲ~ǌ�`gI��RYfɳs����}�ٴ�?���?���37�'���'w��[p�J�C��q�ԁs@{3�� yT�o���ڟ���-8���EB͝3_����Y�(y[�4�?��P�'�b�'ɧ5֤
�qeb����Z�$���� �%��'�ȽÝ'���'R"�~*e�V:q�x��A�;�D� ��E֦9QO<9���?�J>1��?�-Y2{�P� �����;]I��Γ.�\0Γ�?���?M~��4����5��d�7�4"�d��`Y�P���\%�T���DJĄ�>Iö��)9UD'K��1��O۹Dl,M��?���?�3���'�?���?Ѷ�A�d@���tD�@�)�%-��ga���'��'��Z��ɂ�6�DO�V��xU��U�ez��̰,V�&�'�B%^�yb�'E.ꧪ?Y��?�E��&qK�LQ#!8e�	sЉ�KO�6^�,�'�4|�͟�I�?7�E�G	"�#���V�4<�d)�9�Ǟ;���'���'t�	���������U�d�STh�.R��Y4���M�����DVB��S�f��6M�}�t�3V��#}QF�2���*���' l6-�ON�D�O��_M�	��� D�$蔤8.ƌ���|O�p��i�����?��5fj�p��*A(ց�6MF�!���
2
xV��ٴ�?����?A�
;�O��䠟�C07e�T�8�1~O�m�VK%�	96�h�	�;#j�۟(�	��HC�`ܩl���H-��F�]Rt�+�M#��?��xb�'7�|Zc��D�f�B"S�Y�i¶��0�O��B?OH�c:O"���O�D;�t�V8l%9Tj^SM�J���M#��d�On�O$�D�O�d#&O�pu𨂳�q+�<��"���P�GT�$�OB���O��ɡ|*��5����rK�r�MZrѺS�Tq�i^R�'*r�|B�'+��/H�6MU/�|�����?|R�	��D�>Z��Γ�?���?Q��!�~Z�-��<�ա�
���i�Ԡ@i��Jֹi�R�',�	ry"f ���Y�8k�� �`Z��p�b��8Ґ2�Hg�����O�q��.�O����O��d�<q��g��dÌ�s���81��_Z��aƒxb�'��	�d�
"<�;^�(��AE=h� ٻ�Ą�R�\9���̆c���v���a]tX�UK�Qږ�X��_4{�py�Ɓ�F�,�pd�ˈ_5�`�AD�bt��oI���%0L�A�A̕K�n�p�AΔk]B 1�A�N,��Ym]-����8��s�W4R�����G�Y����#z��=�ڲ5E\�1čN3�v�wJ�&q��]�E�u�0��QD�(t`O)���EcңM��}�Q�F�T+�$R��-A^�z�kܪi4d��cH'㨭��a6a�s�ፘ�f�q0��;X*\!��S�C��I�B�r����.}=�v�'2�'���P����$��@���v���eK"a ށ#��#�h��bj�+~&��ư?�=�� �^�Rq)�ƫ>�y��Q�<hB�
f޶<�Ŋ%��Q�g�'f:8�׌G8��tc�7�����';����?y����<!ң�{��H�M��]�g'^�<!�m��<Q8�c�����9!��ۥM#���'��^�G��pm�D�� A�EĚ~���Qc2?���	ݟ<��Yy"�'d�2�t$��I`\��@\�	N�WH�<�,1#1cclr8<O������sʕPp.@#:f�h��ͅ@ٌj�Vr���� 0<O� j�'��i�bktأ�J.3���b!4�ў�F��@.��sĂz �!cD��y��.aD\�Á�*|���,ј�y�+�>y.O
ِKWt}�'��9d���a�@�FԉiRi�.���۟���������S��P���2'��|�RM�m��{aI�Y&��S7�P�'�С�ِ.�r�*%��~��JRe3o7�8��]�:�@�<��ݟ���'�:)� ��6in���S�d����?���ג%	�p0G.U"�p��@��rI<Y4L�.)�́��!p���h��<��J�}��ǟ'?��I͟�ϧbB]3�kS��yc��Zy��Ԣ����z�I��_��S���'�v�T��91
����]�s�"Q:�o�+q,���e��j�֧���ʍ:�2]b�M�*>�@�wDI�V�҄���'�r����f�OB����Hp��� &��Gy�iD"O�� ��x,@���+8]�ɢu቎�HO�S$X�0�Ѯ)em���D�!qk�|�	�$����M;��?a�����O�^��������/�LD��ǈ����D�*9�}⨙�cz�����9T\�UK�nL;�~BIY���>y��ϗa��MY�OǥJ$�1�a�e?�l�۟|��6ekB}�� ��i�Qw��i�FC�I�yT�����א_h� h�H�K|&9a����(x�͒�4z�$Xz�� I��m��ɨZ��!���?Q�����O��Dy>�,�O��؉q%hHpq.�Wy�(�G���n�|Ұ���'.j�&H s�y*FcS}��yr�N�q��ȟ�j�	6*<50�E�dB�M3D�(pǌ�����b����ԑ�6j1D��
�]��zA��dQ�����n� +�}B'Y�Nʈ7m�Ov���|�fa��`���6J�<��� �<i��?���S��L(%f�Qlɧ�I�>6����IBXy���n�cwQ�<y��#tlxD����7������	2�:pk�,���(O�����'���'��\>���?	��#����8�3u�����?E��'�R-/U@��󲀞� CI�Tn�}���M<qf�=T�嘏�����<Q&h�1ћ��'������'���'�pl��h��K
�p��Pc(�����_���T>#<!%%
<�J�j���%� M"@�R| ����O"�1f�	]p)3+T��-Z�"�1c��6�)��T"��?}(�0R�T�0��(�E"D���q-�=H�P3�S�R��Uӆ�=�%���'pb�`v���[��T����C�v�����?�RiҤk�f�'���'C�I��݄�������#Y�$
0�ջ��	4z����� ��g �)��̓�fM0wƘY��O���f�'��Z���Q�`��I�!��E�'B�������=1��B�i-̬�ײ���ȷ
N\�<�GH�\P�SL�J�t��I�5���"|B�bϗK��� (Q$ָ��Ka0�0�fV%mb�')RP���	ϟ$ͧ/U�<��ٟ$����,�0�BGʦ,@,���+(�O<��cX����O���p��$�#-���1.$�O��;0�'?2�O4���z���5d�H�7���y�� 6<Hes���.��ł7M�y�g^ �"qH �
�WXRXʳ����yR�-���Al�xߴ�?����i�|�\�yu�Y�V�AB̚)}c��O��d�O������OHb�ʧ	R�)� �	2\�T��L�!�� Ey-���j��b��VH��X$&�:!��#8b�d:ڧ^rp9��Q�z�2]�pN������8nnb7s�@y��ע�����	<��}ꁛ%�E4��a���k$2�ϓC_Ҙ��?Q�����?���?������9e�N�A�,��Y��d_؟��<��O���I�J�J�c2L�%J�:E.��x�0"<E���:�x,X�$W4��e����ǂ�?���?�����R��U��T�W��&��l��7�y�'�}�c
l*�6��s������ĝ�O aGz�O<� 
��h�	��EЦ!�)�`+B�'��� Mj� ���O2��<���?9�J,�� CT	u��=��l?���"��2�[��<���ԣ&AX�3�K�4*nH�6�����`U��=9&H�)9��)a�%^!�?�b���?���?�gy��'��p�J ���]�8!Y��"]C�0m�l�`[�2�"�R���yy��(���?�'VqCl{��#D);��I��@<� ���A��?���?Q(Oh�$�O��S��>���O*���	}�D9��\./�`��'�bԁ(O�i�*��8�X!͎mE���'<�!P��?)@�ǩr� ���Ą�Q. u�RJ�<�ӧ�8.��!��-_�t �0���O�<Y`
T2dw�Ҧ��n�b@ ��<����S?�j$nZ�����A�d����r�]�A���T�ߗ�yb�'���'�p�X"�'�1O�ӑm.�a�+�H��(�kԖ@<�<1�F�H�O.�܉�.��C?ܪ�#ۮ=���3��$<*R�� 񈩋� τ����J��Y��C䉿|.����(w"�{dMPk���L�;auEQ"��'/ٰ5NǄ�d�I�t6�r�4�?����䧝?���?��eɻ`�Z@�7*@��x�� J=sT|"������I����L�`s��I
V��	�	�B����2NM7�ڝA��,8v��B�n]�z���pc�'���)6�����!ј�dL:e��g�>�S��z����gx�xs7ȕ�Nk1���
9�V8x)���D�d�9%ۗ&��(��@&M���?�'+
���'�r�'��������	�f$�A�ڣ,d"�!pၵw�N�	�u����
^���.R�L���kb�F*O���A��}¦�r�b�#Bi�P�$Qsp���~bK�?��-����G�X�ғ�:v�6h�ȓ�L���
	u� e����9CP���)��<ٵh�2Z�d�BZRUsQ�<Q��M=L1ЄYqg�|O����t�<q���[����B\5uE�E�4�X�<y�Ï*$d�n�- �$���nMQ�<Qǌҗ$`�}�)_(#�V�H�N�<9�+��sh�h]���8�B��M�<�5^g���E�V�
�P�`�o�<iC,�1NH1���%@z��(�d�c�<	� ݸx�\i�ǭàu��i���a�<�f*B��a�͗x)tdF$�]�<�����od�X�Pk6izX��a�Y�<�&�J>Hꑙ����)"@`QO�}�<I��
�s��!��5���Ku�DO�<A�S�?)�J&�;v{\]#SOVL�<� �$��MB�[�X�A�Y�.-����"O 8B��6��,�ÏGp �"O��s�)��K�p�*�N�.ԕ��"O�G�5�8-���	�c�M��"O�A��2�D�[���KP!"O�tj�6e�J�A2n�.U��m��"O�a��.�(s*�
UO��Y�"O����w��� " ,�0�# "O��`^�@6N�Y�-ƕ~��Pj�"O�eb3�
���S,G�GN�|� "O����)Fj�)���R"O`e�Ƌ?�a1�$ϲo�H��S"O�;w�
�K���´鏩�b�g"O.�5�0�"3i�=7�^Mؕ"O❰ �Y����J�|�$��"O�����H+��i�Ip]���6"Ove�|�%�'�XO�*�"O��S�B�"dn�)8&�;(g 	�d"OB����q�΀�v���W�t�"O�-Z���* ���VjJ�"O��#��
�X1��J�xF��"O��S�f-Thd:�)ٯF�)Q`"OX,�i�.M����A�<��u��"OB� p�|q���o3�i3T"O@�)ciUȌ�J�H�y�9"OB��r�H��$U1l�<u"O^u$�m܊���l�{6��Z�"O6���շ�������0�4�U"O�f#и<%V�s%*.�X�"O����B�F�������dm�3"O� �ݔJ�xHG/Ҭk�0da"OfQ����K�X�[���,��DSG"OȨ:sE�8\U���΢}�T�YG"OP�g��
y�TJBmsui "O������h����TZ�l8�"O���G�*����R�E#?0HD�"O��A ��t,���Pn�w9Z�b3"O6�eh_�ߢ�{A2p���rT"O�-[��]�!�'��Z�ȴkG"O�w���l[�����O�P5��"O����)��VŔ����S�=7���'C.��K�0�D�[�H
8�0bg�.�#��!D����h��Dl�m����d��
�@"��5]�h�ᓌU�4Ta�V�by �eڧl� B�I�Dx@9��iPH9+��=%F��
ā&��z��~��\�16�x۱���E��Q#OȂ�y2��(g�`��EV�5a��Ԉ�?�����0?aTj^�`$�;��Bk�2�1l�H�����+l~�	��"�h��	�56xq�����yd�=x����M&?��[b�M���'Cܕi��O����=��	v������uR�L�e��%0�B�	,r4��R.�r
Řu�p^�b�Ab�(#�HA�g��s�\2	^�j*d�AV P�2jX�`�2D����<S�� 0�@�S:M��b<�I��:L���'�J�x�RR��)�'�L�{N��	�'PJ�zT�1z��ڧ�ʸn��I�b���@��+�hYH�E�/
A&I�`
M3U�����I2m"~P
6�d1O��E��Ը�(󉏦#!�ӱx�E�uG�:�j��#HU����z���8e��0�f�
@vq�b\kLB�I�M� #�D�8�1�	%Xb�赀0P��O0C�������H���薨]��Qؐ�E)X'!���/�r��h�[��,��>B��C� *��' � a�����`[���o��U�C�6ⶢ<�%f��Ns�aY���/!�T�G���� �uk !ܔr��\���q/^т��J�B��lk�F�5Y�����hm�uE~2
K�Q2�% w��xUz�e'X>#�!kO"�O�j����$���s����V+.?�ܯ$��rਊ�k�RYi�n�)_��H�@O��l�1k��Gf��HI&LDd�B�Ķ_3V�dF�A�7��h]x�S�$*K5��Ή�� h����=G����i�9*a|Ҭ�����R��ߪY\��`�H�3�*�H��Ar�j5�K>I��Q?�?����H���:W��h�Q�������v� �ǡ�̝2�#;�!$fNꕅ\XP��WN%��O�P�%�s�4�(u�4P�p�%�'�2q:�B����B-�b�R��dU���.�/�X������`CR���Amb� 􄕸=_|���|��e��KżK̢��R�xB�˳K��p?)G�[���!��$đ�'Ypx���#I�2�0�U�#�ZD��NM�OZdk�j�M��ly�.�F��4y1ɖ�"ؐA�-�%
h�uAa�=U��X�k3ړ�DyIa�::�P���L_5q���o�㐆1[�� "�wY^��>I$�M�W�<��7�S:FDl�Y�Fh≸IA� S6.,	묌k�`W��$��%cB����ژ�v4��C��	�Q���3���� ��עp�����|�PZĂ�H=p,�9LO���"�D�O�6]�W�K!=<F��% Y�lBJu���w�<�"Fݍd��Yp�Nn�<\��I6.W<]y�ƃ�Q�,@BX)-�44���`}F1�鉶�	�V�H�~#��蔾Ё��B=98"������P ��;�/�`%�TG�Hj�xC�-QT@����*�=��+��U%��v`_�Zޤ�<�rhO��ޥ�f��3<��ZQJ�I̓MB��Bv,_ $�&��B�M���		$G�BFb�l�إ3�)^��>)n
7D5�x!��h�y�nV�ra�qAPk�� �2 �E�ֻ��<A���7i�x1&2Ba���>L|��'�O:9�f��z��Lɒ��"��5(Q�#�OPLiT�^'GR�yʶ�]-Q�� эC.v�8h��'LO ���)��4u��C�%o��c�l�8GڼEiFO�+_�2�r�� eX04Ɓ/њ�Q��ǅL6��	�8o�=���ս+���e�44|�O��m�[�l1�wn�h|\ܹ����"��y��YrƄw�b����"C��Y�I�e�`MzC'F�\�!0���%9K�>���O��Š�N��[D�!w%&?�~��GM.:kd��A�!?��!���O������C��A���*ZB �e�)
�^�:���Qjҽ*)�j�"�,�xpD)O���" o�'3X�!�9�5ؗC��D����B�*���'J����ITL��E��0�]s��Ͻdq�	peϼ�ē;I�r�'�(C.R�+�r��O����+�|��%��K��R�;��|DxroʼK�<�4��y���*υ�M�O�z�1��V7d��a+6	��?1���d�	�iv����`��x�'����G�2#��xB6j�'l��@ǐ(9�)1栛$#�}�2$@��M��اu7&
��Š�RF����~㢁��@l8��]c��{ԣդ?����O��uU��	���k�_�)�)�(k���dĀ�
 �Q@mˋ>�RC�����a'�,���{�A� �8ET����&�d�J��� �J���i�4[,<�@쟇�V���IC�-I�'�L�0��'Nh�Pr�Z�G\�Ժv����D*c��!��x��Y�+��y�\�9��JɁ�~�O(�e)�!�bl 7$��������h=K�O���"	�&j\�p��ǃ7&$�C�F�j`Ip$�o}"a8*��Uќ'�x�����;���+f���*v�ΝFr��p��(Ģ��ϟBz��0A�hD��`r�*xPp�q���Kބ���ѻk1��@�7Z��D�O�����t��V=��'��٘u�Z�g��̨"�{XfLCI>��Pvl������{r`جj�Pฃm�"�R6zb��ai���3��(d�'�� c�hX�`�f�Jtj8��U�7n������n���C��*�Px�§\u<a�b�Z~y��2���Z�b�qF��c����`D�=L٣	�'b�d��������n�f�^̑A�Z��,9�a1?�'�����ǧ4�5���Oj &��*$
��XC�����QLwx��È���(�UD"��еM��{�J���a�9H�d��#@n����(��-���	Q
�/N��@$���4O��s/�Q��I/G�(`�:�I-C� G�	s�H8�J�0U؜�p @�"6���	�:�U�	ߖC�nE vD[-Ş��J�.�l;p�F$ ǴԄ�I�vmݛ!W{����6)�-I�\��,98"���^�	�nH��"N�v�=���Iq-BX�P�X?�,yɇ�[���x��אdw^d�E�-|����m���~Kr�U������踧��D/�4�λ8�`�ц��:{�����"��A���xO`�CcL�`�b�`�0G��e
 d�l�N26n:[�2����E��8$�p���0{�J��s& Lf.�BA!O��qR�V�s� `0w�
H�8I��흎�����X�0}� �'�芕���9���	�/Q)R�"��J}�ͩ�	�H�}	�����	2'����d��P�'�y4 s�'!�c]"����N�)�z�K%�9U�Y��S�? �q�C��V��z�m�8ub,a$�9<��!� �G]��S�'1j��'E��s�BܻK����/�cw.�Z
�'w�9��WRz~(Z��*P2��J��<a%熠q�� �)S0+4��$��)��y�'J�\\$SeFL� gaz=O��r�&@B?�Ң�Q�����ڼq��i�@�`�<db�9 ���j3�FO2��wB�^�'/$�Q�b�{�Oj��k%,XRf����56+�'����r����������Bl�e	.-<I�'��Ÿ�bRm�g��*r|�Qہ+Y'�%���Ѐt�XC�	;:�%�� ��tQ��;a˅|ϨlC�O[0H�i�%���p>!����	>�pF ��S2�ʄ��u��A8I3�D&�8�D��Ov6-V$���]/l�	����T�ۇ�[�>0!���	���U�'���y �Z)j�J>����{!����&o��M�'9�N�Ӑmʓe�T0*���-�G/��)��B2W�Bi�.��E�P�"�Bޜ�Mf���ы��M���L<Q��F����%�<?Ħ�*ǉ�w8����N�4�1O���#W!bt]�vh�9s��,	r"O�
�&�R�@h��fA�O�n�7�x��̀>�$c�b?ي��$��q�4⇡J	�#!?D�`�Q���.�XM�HHŪG�;D��(�)�[L�Gg\).�����9D�h
�/HRP9sF`;_ ���ek;D��8 +�\��LڄF۶*�����9D��K@o�	2Lhj##M9y�hⷀ8D�dR7���k�5��a���D]it8D��#�J��r���?#Y�<�k7D��R+]!BY���,�0���F#8D���曰J&����P/6�ܠ�(D����_�GhL}�0�P��$YPD&D�a�aV!��i��B 4If�S�F"D�T�)�?s!��zP�˦;LJ���l D��Cƚ.�$1��Huo:��f�?D��Z���<  Y	t+Śl5(�(D��Ⴣ"}X��!g$ZI@�(D�����S�f��1��K�>]#�g&D���e��L���;�k&�d�!K$D����M�$��� ��H_d	��5D��(����\�2����՘|z�j8D���	z��4�fФwt�1��5D��rQ�1@g:m�@�1�&hY�m2D�x;a�4h72��I�J�L��e%D�T�GڿM��lHc,�%FQn(���#D�ifK�7 Y�Q �� M.8��o-D��肬�+j��$(� :RA,�jfa>D�0��H��Rő�ė�,3*�HW�>D�Q%H/k��`�F�I�e��0As�7D���b���
��i�qA4aA� ˥k+D��b�ۺ�(!j�MZr@��Ua)D��P�`ӯ�u:2�)����C&D����!t�v]8������� �%D���
��4DP�F8q�$��H�<yD���*��0"\*/p����Y�<��@ܲf�6�
�������@�<I�ݡ�1"w�N!6�ΐQ�I�|�<�%�n�v�r#�H44H!"Mn�<F&�&.n]c��?n��)�.�t�<��F1
oHg)�=Z}}y�/�|�<���̠1y��%��m����z�<��@�\�d.�5_��D{�\�<�DfP9Y�v�%+��m�����m�<%��06��MiS�U"��P@R �`�<�j�$N�hr�� k q2&HC�<aX�`����@Y��IJ��@�<)ׅQh���cM�h�jM�D�{�<� �D�p�"5�sh�|����"Ot�����h�t�i�&�?b�x�"O�m�ĉX2{�6	��B�J,8�K�"O�ek���Ms�I����/zr,+�"O@���ÍS��l�&�Ėy�X�@v"O��+aa�i��DKD�_"�N�@"O~y�-��0����B�l���"O�hs�d/p�������4��Y��"Ozh3q�حk�b�Ro]+ٲ��@"OH���m c��Ġ�-O�i���#�"O*�:��וt�TIyو%���Y�+D��`,�X���gW�w0��ch3D��@f�Y+hK�᣶ԓS��#+2D��7��o�V)�GN�"v96P-4D� ���un �!I�!6q p2�?D�ԲsB�n���� �֤��	J�d!D��"E� #��C�!J
TV���:D��!˛�lPH9����j��h9D��xa�N�2ɘ�I#E w6�%Ag�1D�TiƎ��U9�Lh�I��#U����<D�l��"^>V�����@1\+�Q��.D� �I^�g���ue���bw&8D�P���)R1���g' �\��\!�)2D��r�L��Iޘ�pu)�`��B�4D�Lâ��5C[���p�Y����b2D�D#5).��`raE�5<��(QJ+D��peǄ��!*����1��*D�4��`��S�!ܔ<���R�-D�@�K�sU"�B��
Q�+\	zS!��i���)H?��!���τ-O!�K38y$��7�к-��`��wF!��ځ}�0����,(j����"eL!��sZ��j��jRܣa`ʹ}Q!�:>�� s����O��y��	lF!�Dߔ77Tѓ0ˈ����@.��C!��[�N�s��^.Mh��vk�3!�Ē>�BA��H%S�Z�H`�.\!�$ؙ#T�4#���d\��i>I!�O�D�^i:�jU�]�^��7��!�8)�FH�a%ЕN����|�!�$F�f�RL�g��<y���sJپ�!�d�"\�l*���d����/��\�!�$5y���P�Ҷp$��u�
S�!��0@0�h!��.�s�̓�Kt!�dԉ(�T@�";��R�l)-d!�DJS"��K׀Z	Fю)Qrɗ�~L!��%%1|��E�`��Io�>H!���TL�Cv� ����ƭ�TX!��;;�.P1,��NL�$��fC!���_~�P
�"�3~6�(��
�?�!�żY��cg��$mQr]�t��US!�d�)xR�3��1ڈQ3� �d*!��Y��X�ĭK�,*�e�q��,!�d �lV�}�ь��Zd��w�x!�$�1N� ����G8%�ݐ�+T�!�$ڶkCdE�U�ç{�ݑeзxg!�d٪.rH困{�l�r�D)
Z!��K�`���jz�t�q��!򤃕b����"h�L[�YcH�;A�!�D@��,��Ƿ%���q��:�!�dǽC���5*˨`ɔ��g�9W�!��1��p�䧄�
�h*d&�b�!�$@��JL�@NA)D�Q�d�r!��[��q��;Jޮ��r#�;[!�� e9�ɪ�X�q`��Z �Y�"O�t�(���� �ɓul�i�"Ob"��'s���і��	l��ұ"O�0Z��W�T�H�E�\NSq�"O^e��l]
�q@Z.>P���"O�<��j��^��xt�ǶzPPE���:�S�@�l�sb̊KT�ʁ��q�B�I<r�4D������@B�-�8�B�Ɂb8N����Y;�:���
]��C�I�_*N0Hd�_��� �|�����>)!̓C��c�S2,�ʼ��%�|��p=1`�S�j94�J�A
 ,�����~�<q���rrl��Fj�dúa �GU�<y��βa�Ԥ`�-�D��Q� �S�<����s�4ŨS+�L�@�0�R�<��)�M
�2p�ʤ`�л�d�<id�˥�h̪�M��GR�����Jz�<�cța�bZj�X�'�4��C�I�#�	�f�θA*܄ ��ܣQ��C�	�s����i_�SŬ�*�.YPO�C�	�3Ȥ�X�CW�9Ή�c،D{�C�	5Rr.���ݾkLb�+�(ęBu�C��	a'�����$4(U��C�6��C�I�W����S��zL��[3c@�+1�C�ɇ;;L��2E�[>� �G�ߞ&�pC�I�w��<��N9�|pi�['j݀B�	#>xz��c��u�B�p��C�=pB�I��}��n�6�2������NB�ɖ@�&Ip1��|�p�""�[	Z�vC�I2N��ŸVG	��>@�4�]0n�DC�I�9�ܱz� ���@A�cA1d>vB�	# �Q�Dj["(:�4��Hd:B�I�`v�A�EK�J�v��w���<'B�'�$`��ǜ�7�`Rfٮ3�<C�ɰq�,ը���^�H���?�>�IN��@�+���^ ��茬v�,�2�<D�D�0�V�h]S�
&�PX/D���b�_�8��-�T) �40��I2D��s�Ѕd6�M��n:S����/D�h a��F�B���O�,���To,D��X��$GEy�C�'q��#R�'D���I�[q��c� �*b͖ya��9D�0zW��&����I�&�8��f)6D�����@#8S�Q nI�~��pj�#0D�8��!
�x��V^���"�C���y"�ѯ�h$a���$; D��G;�O�=�OT�%ғ���{��d����[L^q*�'5��VMN	;�J'�ϊU�D� �'oz�pP��0�X�Q(�-N����'#d���)�!��X�����>����'�^L�$h��uW��j�9$(�E����'xȉ�6��+,��ВL�2�$E��'m����Ǫn.��bH�}.0��'�.�v�˱�d�nА;�.D "O�ѱ5�U Y+��葯Dr�Q�1"On�+��NkfYZ�.F�G=U"O&e[�(�7%0	{1+^b�! "O� *�iL�Kw���"�a��e�R�'��IG�x+�c(f��Yٖ#^86�C� ����"EƆ�#p!���C�ɾ@T��iF _�p�!���M=�C�I#�̸��m��O�h;�/�Bjc���'WD�~�" @	����)�	Hް�*娔g�<��FNW(1;6�ۆy�|��$�<� ��P��/y[PT p � h(�J�"O�l#���'����1Y��q�"O�窆�}DP4�.[8(W���"O�4Iю\7Ba�Ya339��}�"Ot�6f]�@�H��AU�|:l�"Oޥ"f�W��Zl�BK�:^��#�"O(��G�/V���놹�}yP"O���4��@tÅ�_	�����"O��sQ<*�R�Y1��B.�%"OH����IRf2A�>K�:�z�"O�����K?��	��aСJ�"$��"O�A@�w�P`a���b�"O���H-SJ��EJ�\ؒ"O���J�}t�(XQh�-/0��"O�U��	�f%�0ABB�<?R}*��x�E[���O��	C�K�9 � ���K�H%X�'�p��V��Jw x�� �[B �R�"+�eX��@���'}�
	WoA	O:h�ע<D��i�W�NI��B&�_P�`�e�Xh<�UD�>���Z�e΂R�n��R�<�GCԔ�T)u!��Y҄���FK�<��l��f�F���)%�5��BFL�<)�T DgT�d�@�3��}�&�K�<i`lз�@D�c�J�j=��@�@�<Q�ܨSf<PBn��!֬��B�|�<���#4�(�)�.Lz����@JNA�<��G'k����b�#VQӌQe�<��-�ͅ�J������*05pa��c�$R�"ġg���a�T�[��ȓn��I!�/�X"� �`�0����ȓAFбѓ� �N2�b.A֊	�ȓx�V�z�&��C�a�w�ͦ���ȓ2�3��1d6�'�#��ȓ-�.5�-�31ND�@��!�i��	�����MC1cM��Б ��j�1�ȓ#!��3��R�\�+����ޥ���O�Y��Rp AxE�,D���u���^uTI�7E�*�Ҭ���5D����G�8VXQ�'�P +~~�P�%4D����0~o��H�,k2|H�F�3D���t(Y7�l̩Ċ͹�X��Aj6D��6d�'|0|��a���4���5D�졥�^��x�	�LԢ	�*䘓�2D��x�B;Una"0��
����h>D�dX�@��M��-W:k|�M���b�<�0��?���Y�0�r��D�_�O2�B�I��R�zP�V�;Li1cb ��B�aX6�9���.�x��W@HB�ɺ0�@�M+3�����	;B�	,�\����)Oإ�$PD��C�I3�����"�?]�D����ZC�I�hѻ��Ӗyn�ѣ���CA�C�I�f��J��ۋ ���cC��?H��C�ɼWo�hqa!e����Fی��C剌	��p�.؉d����f�
d]!�D��~�D\SGǹ~֬�ehN*hP!�$��0^�� ��hł�
���0P!�1� �`P��W�2��mH�^!�dZ�%��9�f�ܡx�h��i٘�!�	0���-�+�����"K�j�!�D�-"\��AD�t瀠y�$���!�&c�V8�gm܄O�&�xEcٕI�!���_��Y�E_�G�6�CW9I�!�$��t*��4�ӕV��9`��Y/�!�� :��GʜC��X ��<o����"O�4��e��X�x�H�&Rb����"OFX�#Z�"2��U�-3|��"O��r�ϕWl�1��Ȉ�7"O�| ��N�N@��L
X��%"O�	������U��5/���Q�"Oz&jT��ڱ˴�[�M3�:A"O���l�l)pqA�.� �
w"O��A�EɃ	�|q��ޚ^�rl��"O�P1o҄*�2��#�;�LmZ�"OЕh�/S2!�4Bǂ�Qy�,��"OM�*L�1��a�t��Wg|��T"O�̈G��M��c��hU@��"O�P�C`�9����rk�	Bۼ�;�"O�5#G��G�^r��ڮt��'�v�c5��m[)*!�N�f�pP�'0�M0�)\�/Th����,2�z���',z�2DƁ:2-�<:�W!&�ZI��'���I�[78�~��B��%
���'��t��o�4?^�8�)�#�	��'"��Q��ah�jQ'ͭ�bpZ�'���2�W&��<�0'�!7Dc�'w�`�@��SE`9+"��5�A(�'��Q���:k������X:+���'R��p��W	�Ȱ��ʢyrp�K
�'��d��нm[P<�E�ȵi�0{�'�b� &d՞<<X���Kb� ȹ
�'�nm#΋�%xP(c�#��]Z���'��b	�8C�*�KٌT$��;�'ۈ�8�(P���dM׭6�l1��'��k#�]5{#*�@͈�/b����'���*%����ZЃF托�T��	�'�.X*C��r3�]S-�/�a	�'%4U"��')��[֌�2��j�'F �����<��i��U�~t��
�'��Mdhw} �!�Lmq~$	
�'ena�q��,�T���T�nW,�	�'��H��
�75�^d��T.j����']�\�PGA4/U �O�+�)�'�\������~Y(�ڭ%[\�!�'~aP�f�?�RQ:$@���lu��'=|�Y�!< <�C-C�9����'�p$�nK1F��3@Ɖ.�N��'�⼡�I�d���"IS��
�'�vUc'��/DHh<0���[��z�'Vi��@����喂|ԡ��'\�)�#X0�R!C�w���'k��{���3d��T�bE4���'�؀9S��~�Ȱ#��_٠�(�'a&�c�v�`�B<Yx����'���
1l'M� ��Z�V��x�'�����ߏ{�@3�	�k�d��'��;�أs�H�䌒��P����>P�� �d���H�e%*�y2��,�Lʓ���{$�L��!�y�����```蚔u��@k���ycT�	�����f՛��=�e���yBB��J\�U���"r�T�رF��y����|5`�F��n�l�a��7�y���+L̰ܩ���k�ʥ��Y�ya�8-"|�aBHu�⡠'��y��ϓ�P�QDG�; Pu�vI��yBm@$b��W���xQr]�6  ��y�X�/ծ��#�B s���+���y
� v|H�@�!r����Μ%x�TɰP"Oxy#���;��I'E�5���X�"O� 9`��%cc�H����Zq"OL܃bװll��uF%0���1"O.����Ԓ6Z �I�Ĳ���"O�)RK&SMP�{��T2�r`�u"O�`{1N؞#y�D���sx�e3"O�ȠW���I�֠��g\�i�"O��3f,;IjA��.�"5M�ܫ�"O�0��E��X��c�8]7�
"OJ�A���_�2h��(�F1����"O8�ËФ�4ݫ�h�6���1"Ot5��ޕ\��HPH�1����"O*�rA��z7:,������-@�"OHI���˲u:����m�\�"O���c�-0��Dr���?�ȹ��*O�ua��� ��VaͪgN���
�'��K3M�~�|���	�%U�L={
�'2ęf�J.���#B�X�!��'Ҩ�Q��8j���#��.I���'��m�� A-p�e`�έ@C,��'$x �Y4K]��B`Ĉ@m����'R6�AQ`ϊGv0�0�Ií<�vLA�'���vj�C�:�Q��� �%��'���сD( �ޔQ�.��"���'|i1�f��=7�ec�^�}���'/d�j�ĸG�Mxt�Ov�(��'��dD
�8)�t��*��=�����'�j= 1gC�W�3�/[�Z�'���5��Qb:�9����q$!�'�V�qAд!:��;o���
�'[<	y�Hջ"��� BgZ`�!	�'��ݺLM�d�@AwM���ls�'���0	ҧ*�lPfʔ�m��
�'��\��>N��0�� �)����'m	���__0`�ǃ�-����'�~��#�2e�V���( ��'��0��"X3}d�4�$�l��'_xt(�f�0�8���D���'�$���3qQD�iшyb����'��zv�ǁY����!G_'\�^���'���Sf���B�	��I.l�9�'%�����D0H�&�8aA���9�	�'�(:v�G�H��5�4KΠR	�'��� ả=[B������ygZ��	�'p�`�Bϓq��!鳈����8i	�'��ȠѦ�
�� Vg�>�� 
�'�2%R�$F*� �� �T��	�'爤95�B�l�
e[E)U1����'ڤ�t�E� /�aK��4;Nz(�'>����l��C4s�H�=8a( X�'E�D�7
݈$��mz#K�)�x�
�'^p&��}����d!	�AP	�'�"�8r/�<�����
� ��e��'O`���b�-VvAB�-
�^f\��'arȋq�G����Q@�����'�H	�cO8QXZ<Q�߇#s�Y��'�ā����hH{�.��܈
�'������Z�`��p	���n\�� �'��D�Q��2���V%ƣc!Z�y�'�k�&��)�AKU�	.�T��'4T��p`\=9NiCI
�'g*���'��Iw�]�GV813'��.=h,��'����tȞ	2]~Q�특��!Y��� $��0��)
zTȳ�͝;|���1"Ov��'�2�NC�M�|%VyI�"OT�⠨��idX �GA�ػ�"O���T 9���)AN1X@�"O���"���LĈr���E$�Y"Oxū� (g}6����M�2"O���҆L�~����ϛ2��E"O�0�&��(��6M�V�08P�"OZHQ�ect�Qv�ƧW����"O�(s�@N.J�<�����N���(�"O�)ȲO5�T���ÃO���'"O�Qc��6UCɂ��E�5�����"O�����W'�	�L_�~r��7*O�1XEF���P�5�F�}V�X
�'���S���7Gj�+׀ä-y	�'&��U���E��1e��z�ZA��'.X�ѷmȦ�ޅ8�瑭Fa�{	�'?j����Z6t�O�>(�Y:	�'lE�`�R6&�<���90D���'C0h��J��Z0���{�N�9�'U0�+����|�0�k�!
���
�'���тh�%_�%z��U�m~�M�	�'�q˔���UPtq�잏b4�y	�'4�U��+Y+�&�0��B7P�vl�'� ���/�'I��A�"V�,j���'�4�d�HL��T�^�P�'�n��5Jۉ�����DU�T5*�'�f=y��0|�m���1�6���'�X��F��Ӥ��4��,��'�4�6ʁ,!� X��B���pY��'5���'"��G'/^v�A�'}~�x` ��TYN-�d�TS2���'s�<��HQ 	sy����L��	�����qy�,���_�+�f4s��U��y����'D���+"��q)7*_��y�E +d��"t��$.Rx��V�N��y��(��)��Ӷ&HΉ����yB���x��9d�^"$�|�����y�ˍvʴ܂v@��"B���_�yB�CM"�d"j��q	��ɝ�y2��$�
�)���*���y��E)Nݒ��E�
}�ȀO��y�ڶȼA����zf]�P��6�yҎ�4f��8X�/D,E��G����y�Q�4���$�8X`d�0�y@}��@�u�R|�2�M+0�Y��F���C ��,6���@��R �5�ȓ��9ZC�ɣ�%/�U[ m@�"Oؠ�U��m�$!�nC�kwj\�F"O, �������#�`�U��"OƜ��$##�L1IH�`J&�a"O��Y�d�1>�lQ#�Y��α��"O8��Ƙ�!tNu��+�~�f"O��d���;.t��+i	n�<�y��K���i�(*�A&bZ�yB��;%"ܹ�n2�V��J���y��&����$��FqUb˴�yr����X�k��>�j�d��+�y��M��:�*�`��hۄ]P��.�y�-��
_�Hshٮe	.m�&�B�y�H�1ȹ(�홣���*�+�y�h̕pT����};�X
� �5�y�F
{� 	��d̜>PV�;D�X2�yҋ�5H�<�#^N�,"��F��y
� ���/�f���`G"g�ۡ"O��T�f8`h�A	�i:�T"1"O��z�B�57���������2`"O�A�@�4��2���m�t	;&"OH���݌^�~x%�"
q�A��"Ojx�#� ���S�K�*&mE"O����L�w��qj��pK���y2�G�8���jнI�\��� ���#�S�O�А#���u��� cč�+�i!�' ��ⴉ�,	.N��2C�)�5�
�'x@m�S�:S�7��7$e"�"O"�x�cڿ%I�)��W8J-�l�"O�m���*���"$	ӹuG�ԑ"O�UڔE�;87ZA����^�]��"O���� ɀyb�A�V��tO�f!�d��`D��φ2d��i��.�3.!�dͰ;u A���<$߬��q蓩q)!򤙔��!pK8x�,Tq2�ɟ|!������@5my��1C���4y!򤇤�"a�%�V�~w����h! "O2�ū��nV�EȱeيM��I�"O$8��>t��p%R1]���E"O^��`R�2#дS�Fűs�<��A"Or���`%:���$�1,j��`Q"O�U�e� IRt�bѾ2J`�"1"O��RӇ
E��HT��u�&Y��"O�-6*�7,��aB�d�6$r�"O&�#��ěC��i�A�֠2�O�⛲?
���&�)j ��B5��<a���'E�(��ǀ�+�)h��
?�t��M-D��bgfB'<u�y*@�	�U[��B��)D��9�F�,P~A�fM��D���-D������j?.TZBO�c����0D��qA�3,�9�j�a7�Ak�.D��:��A� ��	ǇM22-����'D��Y�M�y��M���G���GI0D�dh�&Cu�������s�pA�N D��ʦ�+�&��eJ=g��ڠ�1D�4`�̜i��K��Z.U����g�+D�؛'�R#'4H���FY�O� �F.D�P�#ă�2�E©�)B���4�*D��To��%�]!�H��A�jh@.D������ivN��ԵVv|E��E1D�����׷o�8;'W�0;B�Fl,D���N���Qg�"��<*��:GI!�3�� 	��^1z��d���э<!�M�FZ" A�gK�����bu�!�� �O�8l[���O���į�b�!��@�<QFDK�L!���HWe!��A�Mxv삵M�xtB�pE"O�B����-4`���1"!���"O�}+��VHm3��ݻ[� �9`"O<��D��6c|�PD#F�'+4���"O�}�p,X�l�E��Q�&lh[�"O�H�UA��VO�ٱ#KŽc�Z,��"O�e�"�DK䫂D�8��ĘW"O���eF��V�!v���p�4"O���fŝcZ6y"��J@`��"Ot��)�	U�"�0)@�U1��ˣ"O��r�i������蒙P��X�e"O��b KH*���QW���s�E""O����eI o/�H�3��)[�a�"O��.�']��u�E��vX�B"OZ����_�j�Y��[�qr�%��'3����O�? ����'ȝK� `����&xhm@�"O�تa���T�*�@�ےiv���"O���ӺyP��q��)lb�h�d"Odً�C��1Ԉ9ԧ��]���"O�1�J_�-�g�"�d8s"O
�x7%���xt�^%1��L g"OT@CWg�N���P��(h�`ⷓ|r�'"^�J�p��;�[�[���!
�'��U�lZK$y�T�PW���p	�'~���/^� �0x�!��!&P`9	�'�@e��=N^�1� B�<���'d*�d�6nN����(5���'8j�*�k
1����M)D����'��E�Ơ^-��i�%�=��H���'x�i{� �_цt�� ��>��'G�q�bԌ�pd��ˆ7H�M�'�>4����;�ސ+�O��0��	�'��{���U��B�ލtc&�	�'�BaVj�*gQ�]� �*s2q��'y��Pa�95)�xI���q�Z�Y�'2Ҹ+Q˝�!|,jࢀo�v%��'��A;D�#O[��Ⴃ[ v����'(L�A�͙,��,��%f�nYH	�'����1��C�0�&l�RT���'���	��vY�0�R��"2U�!�
�'̾2GM/h�ٛ���\�֔�	�'(�@��5X���eۈxp�x	�'ʲ�`���'�lY����Yc,HC�'�����3�� f&��G��-y�'�l�y��ҟA4Z5-ľ:�8�	�'�~$04��WH��D�#�e��'_XuZ4�o��BE#{��'�lX��� r�\]s@�(L�^t��'�:�0��̏f������| �  ���y��
�VA���
�xy&	7���y�"&j���q�؋r����Ʉ�y�/ Zi	���VvCY��yrQ 8�Aa�L�.��%h�y��K>-��!#V,
��z:�O���yBGZE�xT��̵���Bݖ�y�l@�3����S�b�F��ĵ�y�戻-d� �3I�u�ٹDK�+�y��B/��A	���v�f� d	���y��� o��<зjU2sX`���˦�y�@ǚ9��Q���;]Δ�5�B/�y���l��9�u�>7ʶ������y�d�Q��u���>*��]�HϢ�y�ˣ'貹�FE�
(�|�+�M�y�*�).��̋��,T%�� 5O��y��Q�"� �{f��E�z���ۛ�yR.�!7F�i�B
7|$�S����yrɇA�4!��ǵ+���B$��y��[iĝ���J��c�l�4�y⢞9}�J��4�ٮY��1uC��y��ٿP�>��%��A��t�T�N+��'�ў�O� 쑗�$A#���#��=�%��'!���O�j�6,J�>6� ���'+��[eC��YYPB�;d
 }��'��14��x0Ido�E�Xs�'E�مhW�v��]��U�s��1��'t�tK�
̘+��Hbǈgk.��	�'�j�iw�K���
OB�e���'́�o��*9B��d���_֪|��'Oj�i���g(���7nC,`�N����� L��҆
��Ƞ(ڢ2�6]Z"O�(T��
���v�*~�hA"O�����=%�A�P�D��a"O�];%�`�l���^�x��y��"O �b7��$�aJsK���5��It���4	I9� ��$4����g,D��i�'�.�8�*՝I�Nu�#�)D��(�/И����U�+K���(D�0 q*Y,�|��d U�zQ$��@*D�x�eb�` �|�Я�LT��G&D��P�Q�4��dO'��e!`M&D�Hg�W�="͑��޷>5����%��:�	g�'id�#h�7`	ZŎI1C��M��'8D�z&Cy�:���):����'`�Bf�K+x>)3�B�W��`��'���9�E�'G&M��)
/;�^�)�'=�����(��Dj�@P	4���'�8#tI��?��h%O>2j`;�'�2�	��&��h��H$/RZ���Z�x�'iў�O�>� �T�+�����63�5��'`�
� &>���%H�
�'�*��e�Z�<�B��g�hi���	�'��)�#)�)1�fM�l��g�-R	�'�j=;�`�	�J���M;
u�|A�'���ar61tZ�S�"�0�����'@b10S#��%������.�F���'�d� ��L.��|z� �)
bt��'7���kD!�*b4jJ�F ��' �eY'n�$��D���*4/���'��C��f8qY�0��
�'z�U��	��1mRdCC��>)-�!S
�'J��("M@E��f�52�e�'�4P��*l����/<���	�'�@,k E�M4m�i�w��[�'��p�@f��Nh��ゎ�&h�����'I���C���a��h����R�+�')H��Lˏ[[�������Z8�'�,�0s��R_x�Cq�Ȯ42ܭ�'�P��Qkߤ2s0*�)M�%j|���'D�)��N�!1��!��%Ϣ�s���yR/R48n��IRiͿUڴ1h�S�y���(���gҴO>�q)��U��y��-�6���M:O�I�m��y�A����,c��
FsD�X�◗�y���D��1V曹AZۢ���yR�ǉ�6�s�E". ,j�-�:�y�,ݔb6
�l�����'h�م� '�h�h��Q8�r��	�'w����"��d�����X8/�J]�	�'��]{�斓H����R#��uS�q�'ݚI��G� ,� U#�G�p:�K	�'j��  \�V��H��P�~�X�'�d8�wn�4���K�M��%0�'A�����.5\�� J�zT�
�'��F�0�r���F��o��`;�'�vL�%n̈VB�:�y�����'�f��3Nӹ#��ળ/�:?@�
�'��,c�M�e1 Rm�e��i�'(���DO�5��y�B��d�Tp�'��;Q`D�15:1i�+Z�F�̰��'�4�ӄ�]�k0�*Q �A�he(	��?��OJE
0��K�0��� �f�
Q�f"O$�PbhSp�����:�"O��P���hEhuj���"e��X!1"O� J)� R4eM�s��B�Փ�"O�	1��O�t�2�O#A��;�"Or�S`Q�A�xD�f�G�0�Lc"O
�͍5VBt[�)_�%��d"O�sNO�9" ����� �d[�"O�T"�ǌ&:�� �1�8�8�"O`�įC/V?e�C`G']F�9�"O�LA4_�l����F�߳Wހ�v"O�C�Ȇ�l��!�[2T͢1�F"Op1*"�Ł+/�<��S;J����"O$9E C5~�SL�8v^�g�|B�'g�4L���(�'���ekX�5�!��]���JP�M�)�ђK�h�!��."��E��9���{Q)E��!����E�WE>j{r9:s��0Z�!��'9���`D	� ��w�Y<n�!�$\\��*�˂�\�x�#��k�!��Ǖ}G ��a�U�1Sv� ���	�"O���*ޞs�h���c��I�� �"O�d[V�)g��{uB�+�vk'"O�� h��(��h�.Y�7�T�2"O�f�ŕo�d�c5.�R�^ 1a"O1DmKW�ũ0HTP��\��"O@`@�kƀOʢh���2Yu2LH�"Ot ���сM�H� F&�3Ei�'�IO>IIb�*Z3R-�"�! �p=H��>D��sC`ܗ{�V��t��b`}1�;D����)s����/��.�D��B:D���W��3����aX"!'ư���6D�� �A(V<dh� ".6��˓�/D�4I��@=(ψ�@�/��  D�D1q]!ɪ5{3a�
����E<�ֈ���[ET)�� ����g䕰�"O���7�ǿC;hPD�"b"O�ءGԲfL�誔E�'Q��"O��VR��`Mc��ˑ"I��i�"O��	E�b>Rl+TBˮk4�P;"O\و&�V�Hˮ����V�>Px�"O�PHGAD,m�b�� ߉O�fu2"O֔A�6�~t���Q��3"O��a-!m(�H@�@�9:��URe"Oґг(�W���r�͌s�A�p"Oظp�׺SȒK��V�rz�Y""O*��4Έ� r�y��H3ye&01"O)����2r���tŊ[kX�q�"O��i[�_�N�APDA�Gg�aHe"O��@���d��`K R�XtL��"Ol�@���9E`'`W=88��"O�M�֊_�*[���A�''�H��"O6��f�I�+��
/�-D+"0"O�`*�I�q��)�୉&<�t�"O�]��,Y���&2�D4Y�O�)�!��wT���Ґ%�py#W��Oh�=E�T9O|P�׀�N�4c�� %E2�s�"O�-
$$D=\�����̆JCxB�"O0���E����3 Ν#�P�"OVl�E��I}���E.( �\"Ou�Rą�]����L��S�>xc�"O��0���fNusUL�*T��`�"OF�2�NԂm�H����ՎP��	��IW>�����??�H�f��Jgm�3h&D�D��
�Z�$�0b�;��B�M'D�di���0k�����V7���aw�8D��hB)P�-�mה=S�\j`�7D��  �y��V)_�$�h���"�8��4"O� FV�@�4�ƋŔty�@X�"O�9����9T$@�h��çPHXY��'e�O��}��]D8��ue]$z�$ ��:d�ȓ-g"i���>U��"f 4jlx)��QV�5�'ΗRax��ѭ^m�܄ȓtO�$��EP0@�άM�`�ȓU���J�6��!��)��r����ȓ-�I �% *ɤ�JQ�!:��d���5P�'պu���!$^��ȓr���T�H�^Y*�!�M�T*���#A��x��''0ȑ�+U�s����"�ЃcO{y&�t�I�\�ȓ<J��(*�
B�䌉���0�I�ȓX��RP��>|C�,BkU6>�$���x%,�y�Օj,@�FHM65��ȓ;Ȧ�bBCK� �t
6��2Av�y�����u�O�^��Q
�.O��ȓ=����G��$j�� ��#q!��^F��c2�Y�O���{w���m��8�ȓ`���i�8�h�;"@��g� ��M��ёNб~��7Nv�8���(E�U��/E1O(X�lG8�ȓG��TK��BP7� 3 �=2���?���~23�5bހܑrIT�_(�IH�MO�<�s��m���h@%��PQc�M�<���P�J}�/G�-�����TU�<��iM�Gt���pd�qz:4xϕG�<)�½oPA;�
=iИ  RF�<��fR	�V���W;��c�PC�<�֤�/�ܳ£�|�){7�Aw��Byr�OTpx��J2�S�f<.4��'t���4���g �a��m�W�����'�\Q%���cĔ-�T�##��-��'�|4c�OG �ttϔ-��!�'�v4['�ۀL��2p�]�s"�K�'�N�� hV>G���*GB�1R�D�+�'�:UTeD�,(`M��*���HJ>���?!	çn�����jɥVz���h\")0���ȓ�j���OR} RH��A�5U�ل�{)�9���n5 �H�S(P|D{��O��Cn�S_��q��]�D�5��'��T9Tn�86�lE��(8�^��'<��EO�*]Z2|��'Z�Y
�'�%2���5�FL3M4��
�'{>哰�G,;r�)�ꍹ9��@�'=�+ѧ�y TA�I�Sܴ��'��i�M�	n�Xb h��r�"�)�d���F{X] D�~�|�[�×�y�o[�6hh�/x�$�f���y҂��kN�A�p�(k���� )�y��M���Z�c�/j$ܜ3 I8�y��S4"V�)Xt����00�yb� �m( ���d
�o{�lQ'È��y�e�0�V�F�Q<�l�Ƈ���y�A�9�tt��N��b�eCA����y��F�iY -��I�$&3�`���y�;Qq�u�C@^-�vA��h�(�y�΍�!����
�(ujh�'���y�
��>��\����2"���nF
�y�JH&Lδ!�-[�0�l�q��6�y���B���HCc�V�t��4���y�͍>�\��'�~��!dmݣ�y�5�������}b^8j0O�5�y
� �up�c�e얹��-[�?�X˔"O��C��V�t�㦆�]��Q��"O�����>Y�T�(ہ+�z�
""O��j��K�&�T��G��`"OD�u&����&C�*W�F-:�"OFH�0g1,U2��,���Ӡ"O�C������l!`ʇ��:��"O��( ���n�����1��i�"O&��"IA�ı���-[��|y*O�P�$��H��D���/@pQ��'h����])D5lh�����.V6݋�'���BhC<l��x'tJ(�
�'`����ًf��b�.�>d����
�'�yr!��j��L����n�ԁ	�'�Bt��ML���\�@5���"O�)+D���y�d�т+�x�d"O%*�N!9��jw���d�&�P"O��c�͒�MRW��m����"O�B`��#�&P��
���a"O(�j�gׁ:%�8�҄Ťx�(�pr"O0���'�yy��RbdI<|�QP@"O��"k:�BԂDd�Vh�AI�"O���v�I<o�����E1�)iq"O6���̅CT�����]#�[�"O�	#dn�W�4*� �9(��YA"Or��ō�^�4��@G= 8���'2�I.)<N(�!h޶|[��Ed�+�B�ɿT�u��R�H���c�L���C䉧LnI�	[5�M�t#�v/|B�I�|Y�ϓMPha�w��,�\�З'p�'��#;(��V� #]�(�����%{JB�I�+�҈!�Q�y���P�n`�:B�	�b�u���кJ��@�+5qNB�I:L	����$	�k�p��fӃ%�zC䉜)W&�9�K�N>Ku����>C�	��`��d.o��=3c��UqC�I7)�r�pR۬`@�M������=�
ç#��|���D)D�#!gC�q����o�"����� 7��-CƬ�8XJ1��\��Q�qbZT�ԯ^4q����I_�'trq��!�:y��]�-�d^8`�'R�tF�^�	�H�o�"c�f)#�'��cP�Ooy�IEó%�����'aݣ�n\8La��d�C�1��Ъ�'����nK�X\����(#7^r�z����$,�O�!��APh~����eV��:""O|�DV���-�u�ʷqZ���u�'����b�B{uf�p���
9�I�! :D�� e.$�� 8�-��aW�-Hc-<D����ʭnK��1�Ɖ2閱r�l6D�hI`��7}�j<d��$\�P��1�>D�dy��^�\�ăA& {�ꬂ�<D�|j4J�VNL�dѬ''����8D�8+d�U�J�� �D`^���F6�*�Ov�{r!��WT!�C�H��帄�'C�'�az�(�. �=Ѣi����g
��y�ϝ�cL`Dc�!�! I�<��B،�y�Ɨ;_���B�W�f����%���y�k؇#������bd8 ;E����x�¬A6J$B�@W$?��d
a'du!��]Vޤ�C��S�6�h�?a?�r1O�����@,�����k�Y�$A"O�y35+Q*s"p�K])K^(�3"Ov3�ж8=��ID�=�Y�0"O� -ӗ�k�
ٳ�T�H'*AH�'ў"~�@e��l��y����a�5�ը��>��OD��0�d��U!�3�Լ�%�'R1O��h�K��aE��rt*� ~�^d@�"O~Qa���y}\ s�� &\�"O��J`��3N�ɠ���1Z� �C"O(	xMR<.���0l��tDJ��""Od)a�L�������	*sB�\��"O�x��W/ƒ�1cȞ�5F}�`O��$f�8T��m rΒ�0�AA�(,D�����X�h�����[)¥�G.(]��)�b�����N
@N)	��\�A���B���%�v<�uiB�y��5��k�-(ZB\�r"O8('��V%2���g�1H����"O`����(��P�7f��cMb|3"O�𳫈+$�p�
����N��)��|��)��1R��"s� �=��b�F�VF��D.�	0�6x�Š��`�N��$�(B�ɕoS)����v�Z���hc�B��BH(�F]�xjp�����.C䉅��XDn��:����"$%�B�I49x�H᪐8�"Hz�$*�~C�IE|��Z�AU�B��8�D��5�h�OL�l'?��l=;�b�t����w�İh�����R|X�0���~���a�	�M�����@������pJ.�1'U�q�݇�r�uY��bh�#7%��D��������p�»#��\k��5L�=��!�X��#`�`ÔJ�p ��;�T���GA�}�S��$_ �'�ў�|��N�;)h�A���'v}j�y�`�]�	d���O��\���\��<�JD	Ƿc��<�*O�=Y+O�i+�]+K<��I�k*.��e�'�a~��M�U�LU"��υ3'��������yR3LX���g�,2��B�yBeG�cXꀨ�n)�u�ŕ��yrg��:4<D��P�:M&b�y��[#��U��C,c�H2������'�azR	Nmr����cy��(�l����>)�OnlS
ڿ]� g+Ғ1p���3"O��j��Fu~�5�+W�ns
�q�"O�\aU(O[���٧O�T��"O��y DY�G*&)�%��e�2 �`�|B�)�Ӕe�� ���("W��+�o�4!OC䉺O24 ����`i�ɲN��Op��hO`�	� �j\P3o�f���F�Y��B�	�oޜ��c�P$T�#@��$B�I1^�PQj�; ���ŧ�	FB�I;Q�tEڇ-�#qM�|��`�B�C�I�V�$����}��Xc�����C�	�2�轺�A�~l̑��ZjC�	>�F��r�[�e�r��r�M-��?����B�T�� Ң9�v�x�F�(!��ّ�z��&L�}�Q���h5!��3y1�Q���hf�8 �`,!�ΡZ�lᓢa��D���v!�Č�	2ZA�g��S��P�n��B	!�$�]Ӟir�˙H4�R�.��'�!�D�"{L$̳3cQ6N)��4�ƚH��O��=���}1ܑc���*��Q'���p�!�ă?-F��P������M7^�ў؆��$`
q$�)��i1D�HC�	� H�<�VO�-���7u��B�	
Qx�e5iґ=������G6t��B�)� �EI6\�p�	8eQ6��%� "O��i��z?��1� j���"O�������Z@t"]#v>���"O�M6L :O���4��,j��x�"O�1
v+[+udM1��(4�"O�\���ݚC&��"��u�T"O4x �D�*"�����K٨�7"O� �s�A< (��6�I� bdL�"O:9;'I )��<`ѡ��b�p��"O��KSǑ4#qj�iTA
�x�"O�,�<Q�t��� �[	�!�"O��ae!��DrX��A���@�JA#&"O�1jV� �Fu�S�*��M�"O�䳧`�����S5/�<�r0"O�u�@f �T"5%��Zx"O"q��������*�?�xa"O��ƣK�b�^U�"���挭@5"O.I�W�A���3���-u2�9"O�|鐥�-F�
�2J�("�ҳ"O.u9vd�r/8X�h�0m��Z�"OT��� �s�B�C5�JQ|<��"Oh��v����ÁZϸ9�a1D���bǜ�q�M �k���7H1D�`��l�
vTPA���c�.9��;D���H��i�$`��	U"�H��,D��i���&p~đ�!�F�G�ð�0D�p�M0i�6�г+�-Z�,��&�,D�؁�d��c�@����p� �t�,D������%� �PЧ@o����� D�,;�,�B8��X����e)�k0D���b-��a�K ?Eh�jci2D��CFIT�e� �bA��ߞa�	/D��@^r�$�!�ߩ]�N��n�zj!��M�Y,�t�%レG�f�1��U��!�d�aLy�a��yq,��`+ �E�!���v���U�w�Ҹ��O�J!���i���q�H���L�B�!���X�4R�>�������bq!��5s5���Di/nn\ܣEk[,VY!��?�~��D&
/j�Z�cC �!�DÛQX>�J��`&9�B�9�!�K8�lt+憃��hr!HL�!�d;����a��!�Z�!0M�Q!��w�F�z��;u����A� 6!�\!c�Y��<
��ȳ�B�wE!�ĭz),��T.�)*2eR`NZp.!���2/D�e���%��l���ΧH!�M
�<
�m@�g����70�!��xi:|�s�Q�,�,��#�2`�!���7�XH�����h�aBT��!���b����"R=F�Ht9���&k�!�$L:�e��D��9#���u�!���pIy����y��F�@�!�d+9�F�i'���u ���	�|!�^=�l�f��Jbh���^!�d�G�f�%��Xn�b�(Y!��?(�����Z3i�%��!ۚ@T!��E� �|��uf�2T�^h"�i�oL!��L�*�[&�ַN����0	�h>!� M,�,�DG�CT�UL�`\!�F�V�&��QN��\<����U62O!򤊋^�.-��J^ r&�A��m)!�E78�&d�U-��^��Xx�K�j�!��
F������?
Y��#�Q�!�� v|s���Z�:�!  vf	8�"OUcf�R�]��@�!u��"O.l�p̃�_�Ta2����
�H�r�"Oҡ���X
 -fL8�)4RR$�a�"O�I@geY�>X�B)�3R0q� "O��a$�ͥE$����^Sl(3�"O�����,QS���M� v7�M�"O��i��_�W��#b��(t�"O��r�B�y�R��l�3�b媱"O28�mY�
$�3ՄY���b�"O�HIEi�R3@��.��@��"O�HH��H՞ W�D�"O(�;�"O&l�G���@d��,F'(��	A�"Od��V�̰q˴��&
G	�4Q""Oд�vN^�mR�ږ��(���"O�)P��/����`�҂]Q�"O 1�f��9��\��f��z"OR������)H`i�D��^d�Q�C"O.��֛���j�d�;E��G"O�+�!��'��`����4���6"OP�St#�)e4̴j���z,�{4"O��RB���;R��끁F3ڝI�"O��)����\c������	B"Ox�e��V�BcGjD'(�Q�g"O܁��A�6>���٥�% <ٱg"O�-�f��d;�E[�'B1m �Ȩ�"O����@�2�,���eG��@�"O�BbVq��1� Z\6%"O�h%�ÍB�d�z��ۼE�D<[P"Oĩy���vN��D��B�f= �"O�0RrH�$%�	q�B<�L�9"O&�k�E�"�0HS�F�`�\�u"Oؙ����έK "�g���{�"O�����V��5����?@w �i�"O6E�K��pN\�� #*�85
1"O���B��\���.��e>����"O ��苨O�0ԇJ�% qC"O,��a�mkBU�g�#8����"Of�@�'�ojF(a�]0Ot�0�"O6`H2HD�G���Ԯ��q ��"O�P:& K�{�R]a�OD"Y�><��"Oځ�5F	Kd�Pp/O�L�TL)�"O���gEI>�((���z\��"O@��썵K�(�tϒ�%��01F"O��s��/��ŋTę�y⁁�"O4Њ@鈦"�.���"��	N%b"O�����Y�jhnUzр5p	�a"O��c���5>`�	@ ֜W�f�PR"Oi�Ο���t����!����"O� �JD6�<aQ�R>0�^`��"O&H	׸>m��2g��;��;%"O� � ��@�=���6x�6<�w"O�����0P�ek��P�^�vĈ�"O�J�<oJ$��wMįD����"Ot��  9.7@��)^!锑��"OXDZ k=x����ŇS#4�;"O�I{�FМ( �yW�7�li�"O.��R��TZ8�g���.���"OzpK�$?�����F"g	mH�"OZ���&Ҕ.`9�Ub�0.W�]i"O�� �	ûb��ˑ!ؾ)A��z"O��kֈK�e�����mC2"O���瓕/b���%̶F
D���"O��VK�?!P�qBs˘(i�郆"O�  �"���D$���Z!}j�djC"OܔR�L?� 0���_M�b@"O�l��\eҩ�&��N��Ҁ"O`�y�Ǉ�C
� �d��25��"Oёrcѿ�r`*�ݣ�Q;�"O=���[!Q���36�� \쁔"O,�٦��<�^wF��\$ �"O6��O$|T����O3#�:��`"OfT�0��%X��� ��ޑ&��h`p"O.��1@��,��I����GCh��"O�UY�H�0����bA�R*J���"O�����(;V@:�Cȏ~$P��"Ol��)��
����`��<��e"O:d�Cّ&����-НcfL0�"Op5@@cN�LZ����K܂=8�s�"O��;6B&W4b�A�:B}�"O|��f�#q��[C�L6P �@"O���U7t����D[DT�BS"O~I��[oJ�*��;nh9 "O��{�iS��T)3B�>[�,��"O�� ��N&�t�u��v�=�b"O�-	 �K;U�F���1��ٗ"O$a� A)0#��[�oY�3���"O��h���c���ծ=g��|J�"O�����I������
Q���Q�"Oh*�,����	t̿�( H�"O�4�2�N-.Y�EVr�`��"O�y��L���Ѣ�%A3}ƶQs"O�ܠP�B}Ȅ��D�v��"Oڈ�1#�#����`��<+�"Ox��%Cݩq���B�W�HN���"O�I���)w2���	Z� H�P�"Ol�H�Iđ%�8��F��DE��q�"O�u9�/ؘj�HV��#D�2W%!��V�������+��d[W#˪,8!��X~Z:��	�7�pYZ��׾N5!�M�O^����Y�O�Vd	�˸
?!�䒋_p���䇾3����e'�TN!���9�f]���M�z��$�d��x_!�DF,{��}h&���A�y8����Y!�צqJnH�B��ʪ���*�6�!�DL�����$]�&�(Q�T"cr!���* (Y؇kƕ*X>�+��2!��`Yt�J2V)Y�!3�g\�!�Dp�2�iS�U�V�<H���ȓfa��Xu�R30�ʐ�3�ş|�l��8���ؠ!�/<��j�OD�����"8DPh�*�
R����׀��%�ȓ��(���|d"�!��R�5V��ȓ�����T{�Ɲ�p�O�:�هȓ ������A�I�%�Ł(.�m�ȓ]������V�QJ�Y�fO]<E�ȓR�.��D�!Q�̈���9W��a��`sX)�e�C6^R,±,��8=����	���(��ˬN��Qw�8H�����]q�#��8Z���.VP�E�ȓ&�B%���\?8��sg#�$U�@ ��2.��r�IJ�m�~�z�h�&]�B��ذLi�.���2fL�9+,�C�I	k� ���Q�4	�vQR��C�I����$��.W�Ɂ�#ƾC�Iy-­k�.�7��$1ӊ͏lO����T�q��ԥ*����)��r�^צ����՜!.4���� �MqH3D�� �!zR,�5$��\!$�,{��t��'������.)��D�l]V� ��\�f-�ȓ&���!m@�&�5P�х�5	��S�
a�~���)r���^�h<� F�l�$$PjH�l,h���ɘ�H��	'0����1+�?f���#�ќq��C䉱?[R��4�]v�:�5/��F��C�e���r6@�Q�j�e� kN��d�1��jX�İ�����H8Ʈ@#=R����j��棛�w	�Pn��t�=�������S�;�H�V�ߟ���qn��yRIA>�.�b�l©[1�x�'�W��yª�|����@h�l9��>�y��U�l������b1z��E��y�Eɳ�x c��˘g�,RB��'ў���ѐg�=7��)�2	�5biKv"OI���P�"�P�S�i�.�H<����I�R���s��6t����w�4*w!��J�!46=��� |D�5B���5eBqO���$�
MI��bD��?��0��3B�y��xR�Oഩ/S�<ׂ\£N�p����"O�q�_�H����Q:[-���"O���'���ѩ#
Ԑq����ύp�<���αf#,�#��Ҳ����e�r��0=9��:��M�ӃL�xp�T�&iCY�<aP�]=H��qB�§�͂���\�<Q��=k�~ڃ��"ss�}�S�]�<	�OLE|q�c� g�%J�o�n�'��y�擊>�� -ܯ!��z3͖5�y�&�gy�}���D�	7��c����~��'�f�����%Q�� �,$�Щ	���1��K�ӌ{Y�4J����z���Z��B�	�eq%BI�1yb�e<�B�I&5��D�BQ� ˆ$ҴX�}!���~�t���+A�6�s-/G��O��hO�B�����'�����S"͝�t!򄘚H�~y���_�Sd��
<f!��D>3�:93f�$o?0����[EJ!�U�J�>�c �M�12�4����55��]�i��}��e�_�<��D¬"�`B�	/,��B��@w�t�wlK��t��$WZ��;�����jA��`�i��*A�1�ȓA���r� ��/�A鴮�/PL%�����ɂN�j�'�D$[ӈ�)��97-P�<:��
�'����SŘ�v�CA�d��dJ�'A�,ݶT�#"�+P�|8�F��|y(C�	�T"ny��Ϫ4)fLz�cL9�B�Ip*�T��
�	]�Ī��uW&B�'P,�0�c���"MQ�%[2��#<щ��?�5G�+p&��DJ�1:��&�<D��0a�=���K]4b��6�6D�dX��ϕj���1A�@
�EH��>��������BQ�Dd+�$�U_���c؟0� ��#����kC��Q�,�����<�eeu�(�h��A��-�c�4g+ =�å�OB���C����t���
fis'cΟ�T�>�'�7�'.��ƍ���h�5Wf@����\qbS���|K�KÒp��Dx��)j�LȒL����#�;A���H�K�H�<�al�:v#�������jsةH�*�|�<qAN�0F�	K	�%�A��d+T�$xC+ �~L�*΂!!� �A(9|O�b��r2�E,�V����%z�h Ph#D���V�$�;�e�|s�� g�;��L���g�? �,8���rwR4��յLD��pw"Ol�ӂ�ƖP�<\��e���68'�>(O�����Y�PR���t��Ycg�Ȳ@(uH�>D���-ߑHЄ�ر�z]Z��3%b�8Cቇz� ���Z�47BЮ�J
����'k��).�����:c'^�6g�M �O(��$�:jhX�S!���$蘖Ȍ�&�O�㟰�����17�=��S#c8%2,	!��K�ެ7)��~�b�	t'�)��O���'�)�ɋ-e>�ib��Ǝ$��B�Y��!�D���};C@Wh�Na*��_�!� q�D :�Ȁo�Ȁ��V�z�!��Q�t�ư��ܑ0#v�Y�L�{���Xx�����)|��b �=4��U�/!�O�ʓA�|� �$-(x�ra\,.YJ<�ȓAN��"��ܻw`z�#g��.�p��ȓ	�(�A��we
�ͅ�Zs(�͓��?a2	2-���3��J�_��ٵ�E٦1G{���i�ƕ�`��_�M��`�+���X���6��h�z�G��7R,���r ���?ѧH�)2T���'��w[���R`�<Y�%fs2�B�Bw.��qF�a�<ɂ��"?�J@���'Ny�Ec��~R�i���)���I�X6NU����&G	�n�x��/�O�ʓe�n�Xq�3	s���fW
0>��m���t�?�g��?1G�޻<ج���סY��4[�<y1O��,��P�љYp@9A�V�<���2v�T�e����HçI
HX�ܐ&\�d� Ȟ�d3����J�f�$��7��<�S�B���
P�N#(9�LA���r���=����T��D\<�`�U/rs��r�F���'�z����q��i��-7�xᓢ��(�M�3;}��O?�|&�pK�b�ڒ��Y4�|�Q�*\Oxb�4"&�JAn갹�Ɵ�,�����&D���CFAe���4��t�Be D�����s��ź��д90V� �1D��+hl�@�y�L�??���`C0D��0�A�%d�^u#!��
�x��4D���R%�%��e/	�h��D��!����	3�!;`��T_�y@�d�%a#!�$/`~A��h��3F���c�n"!�D��tF8�37�4,���a�0!�D�8N4	1� �` ����_��!��A/sO*�����p|\�C���K�!�ԇ5�&Q�%��'5�P� W���!���d��m�qD�9���J�[�!�$@�=�l�Q�kL�wf<<"�I�#�!�D�h���樕tv��Tg@�@�!�D���І\g�,�!�c!��r�l�bEH�T�> 0��R!�dȬ{��s���q�.�F˝5n!��+1C��`&�Bz�.8;ď�7Y!��05j9��j��[�Z��V쎹O!��?5Ԛ�h�+���U���f/!�D�a�lq����Pw��"�؅h!�d�*e`�B���~f8Y`7n�u�!�DX�RΨL��7,뚐�tπ7 �!�Ϗ" �������Y�g�9�!�92�:DJ�j�d��1�7	�L�!�d�Hڤ b�E�+	��4j�
� i�!�Ӿf��
7��('#�k$DE�!�D�,����%�&#�ek���5n!��2Ch�U`2�Y�B@�
:S!��ݴ�>H�Wcߘ�D#u���!�� Z������.��P���@tL��"O����jU�,�3f��2>�
�"O��h����T�M�""��jb8:�"O�Dc��^6�	"����c��$��"O��Х@֋l6 ���5{Bh-�"O�TsAgY
p0I�Ϗq֦Д"OX�r�G�0928�5o j�fX(#"O�d�7�ʠ,�UӦC, ��T �"O���ܦVQ�h5Cŗ%p~A[�"Oܘ�W�(.P�h($#�SYV�H�"O���g���$�tȆ�͟D�,x�"OZ=c��;*Jh�� �7;�*D"Ox�k�*�/\Mb#F6��X�"Or%pqΙ4�#�Νm% ���'���b�@tѴ�*�H�0�9�s#֘���J�'3z��7H�z�q��Y�=�R��'!ꥣ��(~��Bn��OO,8��'���SaH�,\�rM)>����'���R�L�5�V$��J3"�u��'�xMo��V��);7@�*M ��c!"O�h�m�)4�j���;G���"O@�Cte��'L"�bvN�2�䁥"O�h�fMG�Y�F�y�Æb�P
�"OD�:��dc�p���ʁE��p S"O�|� O�]�8L²�\�}�z<��"O�T"A�
�f�Y��ץ<�H��"OJ�:�!j�XDR��PRj�#�"O��I@�X<�䭳X�/L��"Ol���+���Te�$v4l���"O�jt쏙z��e��
��n`�Y�"Ol(1��H#��R�G��R v��"OX`д�]�b����S,r��\["O�����M�B��a#���f��2"O����P��q*fHV�_=p!3�"OjA2 �%�>Q	��s���"O�ts3�G<g6�PgM��#�~�R"OXt���-e%#q�ep��f"O�}	����-���5O	�c4"O6!H �ݭl-HHT�N�l
�|��"O-�E��0.E !"�^1J�
ۧ"Od5���ٽP�y)0�X+t�X=[�"O��RT�ڋ&T@PR�Ό$��<�C"OF1j��Э3pzQ��NH�|���D"O���u��@\!t�J�PR�J"O�[£P K�4��tm�;�l��"O*eI3��W�������4db��"O��@��1O�#��B�J�4`R5"O����HR=6R���%�@�tJ0"O�eS�c�:��e��ǖ8���-�y�䆓"dq�堞:*28��a*�yR$��n�8�B�B�.*4�����/�y�&}�Q��%�'Lc�<�fN��yBNߨF�����u�CM)�y��& :Y+��90�Xv��y"��s���ӫ��~-RVHV��y�×
b9��	�H͚}�l���U��yB�:�d��ҫ�.g(es�
��y�O�L
�ג&���"�(�y��F�|�V�s�*�6��|���3�y�"M$�!y$��W���EC��y"fF4E΅2sdJXQF�ѷ����y"C�'�I���"W$p�*"(�y����`�D���Ʌ�Hʔ!����y�LS�#���Q��T�A�f�*�K�-�y
� �%RF�)�t��'�!S�^��"O�<��A�<�Vd�F�#a��<3�"O���R�&'F��`Ƃ������"O U��H�V���pe�!h�l\;S"O
�Aޅ�|��
O25B��"O�)H���+�`���k�)�""O��'듒,S���W �l^ ��"O|@$����1��	LO�( "O>��!��+U|l!�q�V,��B"O�q�F�q�*�J$�,`�y�F"Op�Ԯ�+`k�3%�L���"OXȁ�O����)��
B�z��v"O�qb�����7L��ڞ� "O�LfCw1H���E�d�z�"O���'b��S�
�׃rh��
E"O�Mc��G��QIe�Q�wn��G"O�d���
y���0�V�d�V��"O2� ���$�
1Сۋ7���Ä"O�����w�r�!@]u� ò"OL�*���mP<�� \:+�PA�"O��{�{#d�`�bĊ0���"Oz�Sqʞ"�>�B" ��q�4�SB"O�(��#�!:�����������P�>���]�0���?�X���0ܼݫ oٶ:�hCR�5D�0*#NԪ}G@��R�V�yf�A�$Pc�	�xb�i�d0�3��\�(�r�*q~\�{F�D�V��ę{JPU�� -��XYS)��޺��$��'0B�x��7����Ĉ�	�0���%���xP�X���BPkܐ(q
�m�3O0ɑI~Z�<j����N|RܡB�4D��*�Mf�!��a�l��I!&�/`�� �^9x���b��?ك�2_ě����\<���y5^Р��գ�y�ߪF�|�#D�)v0B���P��z��=G~��R'�S"R��@)� �+E�t�'�D9��GT�(����rYZ���n�;&Vv�9�[����pR� �V�8}��ڲ"�7P�Ҵ�q�F���×!I-.-�tM�(S��S����c��hN�Z��J����,��ct����&!<Ĵ��06��Or�Ƞ�@��j�}Q@_�H�X#�'�TM[����M��	<~�6��/J�I�T�!T�]�&����W�=M����d�D�A���`L(�!p�ni�D�>m�nXPŅ�-1;2�� O��<�l���"O��R�c��6h,�Y (�n����Hn�~�RF9�A&��v���UjF�)`��'�-�ݏF��-[�&� !V�����#{�Y��ɞ( %���Y�C�������	v�`�SBB�`I !�R@	o>�\Ƞg�?".��Ox$����'�\�a�Ē=ehJx�rCc�]���D�I�ңj'~�����I\9�fQq���"h�$�(��"2��Ċ2v�i˥F8�0=ɱ �"H��p�V��bX�U�HT:	 ��)N�l2�d֥�<��h��bLK;��r��� E����d��D2��$�l�9�'���jE�P�[�!])z�R��4�Ra9�H�vO4�#E/���0�;P���~���x�V�'Gj,�
�� �u��M��C�9/ڐ��	6y�h��&n�4����*;ֈ��I�8,�W�_�A���3�H�0� M�j�5�'�3}ҁ/@�J�P�H�ES���$�фҸ'_TQ����(Cv"J��D�q��j6×�7��H��C�)s�)gɟ�e;h�*�/���>a�D��}=��
��e � ��̃N
l�Wc�*C���I&@�=�,�O��r��<�<��'�Rj珌�>�$�X�L�uߪ�
�'�\���+����d�>��m˄]�T�����+
L���+ڤ��'��i��W���t��qCD�0��2Q+������<9��F3R,�ɐ!b�wL� '��5;�YѵN�I���T�[`�y�S�8}�	�!���v��L�B['\xPc�ײCS�� ����CP�����)V��dxf�7%�p!3L~2f�%=֢��%ťFLN�b��@rp��m�]FT����n��yss�Cg�P�ƙ�ad:x��J�1+.����h�06V>��@�oX�yvP�`q�H�_��[e�M?8K���5�,4��@L2ZA �C�@Qh�丸�bH��<�dA=3�����[(�h�H>��KO
Y-�`ͧ����B5�~��3�E����	�4�t�����C��3P��-E�A��
�i�Tn=\$�2/�IK��s�I)�dW0��%����LYF��B��@�D����2�S*�r:�CP��t�	K�Z,��u�� ��TY]D���d
4uC�I,� H̠�)޽=:�0 ��AI�ٓ�\���;q�R=xt��A?@؈�^=��	)?�Ҁ�*0F�9#�G�~x��g��]8���&L���qP��l��k�b�L!s��҄=�td��O6>�<9�0r>m�C�G,b�x"�K�	`�x��;B'>�!#���	t�^Tp�B�-7>�	>� ��0F��\bh��mn�,Y�"zkN��un�?�M��
O��3#��v��X!�Vs�H�@bǏ�1 ��t��!��}a�q�Nۚ�?90ΗD��݁`zu0�o=rH�i�F��A��C��0
�L���k_�x:4�6L��(���IfI�=��]�׃@�h�P�I�e�X��c+�z8�gy��
���X3�f�*DH$� �p<�B�M&J�q�@a1?Q�U�G&pZ��'E�"@�3V��$��Al�`J����<�c�G0%'�ԡ��נS?��97`^Q�dU���ݞw�%��"�jƺ>��3���`����-��Y�5;�o�3f��
�'�X%�)�:o�vXr��.�[�(�2��9_ C��*f8�rv�(Xv�}ޱC+�	�Rh��Z�c�N@S�`'$��GI^�	��`���6=�����b���!�`�
��I�+% �#d�Ӝ��gy2(C6"����W5�4Ճ`�C���<����4�6OhIQs~B���Ϗ=6��G�7��0�����a|A�|a��[�5w���:`nY��p=)gmݷ3� �s���x��]a4.L�\ɜ�bG�ر]��:'�G�Ɛx���>]�1 c�A)�%����8��'���c�}��dy� �A�q��T�"�.)�F5s��:n�\�"O�Y����0��K�G�L���Cܴ�U)�(�0Gx���Ծi`p"}�'K����JV�m���`��\w��a	�'Č��ᄩhn���A�U�ܝ�C�0@�����Jy 5ݨ�0<!ǄR� �8�DD�m��a
�p���#�l�$~�Vhkv�L�L�iK%��P�+�L:q��	�I�!�¼p�X�;��E�^-���@�/�I�J69j���a�L��o�*S���4�c�'�����w�j`� �;]�X��8E*	(��:k�~���D]:?��pӓD�e���J8OԹ��H�v�/4z��c�O�E�r��o�h����%���:��'���2fM
�-H�|Ir$�gg�	���$"�'@�YR�Ͱ5Ί!3ц�&&��Ĉ-x��
�!	6ԍ���^N�Q�0��'��e�� sA\�7�M��H�.�qӗlf]~�`�<���*Y6|�!�D_�>ε��A*{_�a�'B�[���E�TJ雲�Ҽ2l����؞�PDX�`�}ܧ~����ՂP768L}�U@�,��̅�)�f�Z5�\.=xِ`�(E��d�R�(W�����a�;�*�+�W��C�tO�� hm���7��%	*8;��M����� 	�t��VB�5�b�uP�7����i"~p@�jF�Y�a|�ӿU 8i�eb�j��$�U�ւ��O<�k��$\,2`�f�-��V�jk@$���TY̪��F돮t
!�O1/�L+
0eBj���J�DJ8ZW�5`�КfnF�S�O�P�2S�^�w�P7L(iR����'[�z,�5%�	d��c���z��>&H^�E��M�՞��}"
фu�"XaQ*ʗ4�$	�U�]���?1JQ�t�8�x���(ZNv\�UE�1V����Ƀ�x"oҏ���b4`����ؓn��y� "��sd���i�@�C��%�yRDB/\�p L���d�2�M7�y"�֊,�� ��S2ʞ(�H�y+ǜO���"fC�$�hV�D	�y�)�l"t��P�J�
�f�B�7�y��I�^1x����^2n�Å/A�y2��u<��d�C����å@F��yb��	*����)K $I��� �y�`I��TcR��5���A���y�Ȱ-
��Vb�+�\Z���;�y���R	9f��%�8�4a��y"/���g�6��`��ES�y�y�.q����!����y��M��q�'l��|��h��OT��y��5:��M)1N�D;r�����y��[�@x�H9lwD�	&�yr���9�Uae���
�*\��j� �y"�E���*��@w�|*�:�y
� 2�c�:,�҃㋗�\�r"Odr� �9̤�fh!wFE�"O0���=��S�G�)}P)��"O��@D�?�*�3�I�	�)��"O�	੏� �TX�&�;��U�"O�A#T&��zW��QK
C���%"Ot�9�*�8�N�aS
�%kh�"O�1����z��Xg	��*�,L�"Oب0��10T�Jg���6"O,�S���S �Y�%��"��i�t"O����J^�la!?p�РR"O����j�}|а�6�s�<@"O��rc�ɜ!�*d��G��z8"O4M����[3�U�' ����p"O��sA�XL����P�W`~р�"OF��p틀A���Go�p��8g"Of��1+�JCt���Y8=袍�E"O4؁��Ll�4�v>d�;6"OZ�׆X+l����L9�'"OQ�v� 3������~���"O��pC�����7����"OԄ�P�.g<�`��Z^�pH�"O�d�ŊXP���T���=����"O,|;Ac�q�i��bK>�*�g"O����㏷||�p�!�2c�r"O ���A�>?��qvCN�z��tK�"O�h92�d��d�!_t@L�!"O��;�G*0t���B�Au���U"O�XU�Ur�j2G�]@\)��"O 1�qj�-x�h�H10!6�"Op���M]�y��8q&DR,��!"O��'j4�ZbD�#D���"O��C�ֶ&t�e��l�T<�"O��e�L�.��]�&)�~�Q1�"O��M�=$v�{�ʕ4��x�"OB��m�#
����T)2�|p��"O|i��!�X��qʏ�/��Y�"O��* -��a�Ȅ� ��*F���D"Oe��M9-±�e���n��8KU"OHX�򥉃x��p�3���rQ"O��9��-Q���[���sTI��"O��TJVN���2CO�0�Ե "O��R�KE4�>�C��T� M��"O0����Xpӡ�v��AX`"O�����݁�N��%@�b��Ё�"O8)��N4o}���$ݑ?w��)�"O$�qL�L�dl�c�rVx�`"O��r&@�%_���p�hM�`�5"O�ڣ�C6 FLPW�[	cO��c"O����b�䄸�� ڐ5b�i"O����*�ms
��	�>�N��"O0����"~=.�k�	0^�mpU"O����"L<��ς�U7�@��"O���w͕7o�9 �N�#�ظg"O �w��� �����G�Z)f�*�"O����lq:.lc$��47���@"OxU`T���l��(��H�o%���"O(=	D,�4S��X�+�3$%�d2�"Ol8��`Ǿ`�v��Ζ� ��"O��Z3�.50��t�@!2%�A��"Oڈ�Q
R4K���c��/4iC"O� �T��A���P�O	�2nh�7"O^y��̌�6=0(Sv��3C
� �"O�D�Dn٫YK��b��4�P%�y
� &���Rl�>��䅹,P0�"O�$z�O�s������O���["O`��q(	m0<��P+��l��"O�l�4(�y�fxᡇ!k�^��"O���C�Sc���7�;p���p"O��fŒ�9ʕ��F����P0"OJL�cǣ?�V�9�d�>D���k"O�0��ىXr��sŃ��!���p�"O��@%IW�n�0C��A�'@;"O�a#���!���!MIdk$@a�"O$��E��a4������@"O�	�g׺l:��C���7"Ot�4
���&Զ?Ӯ`�A"O��BRK��b+�h�j��O����"O�гD��2X�, �KƼ$O,�7"O���)�/s���ԅ��d���"O~��ej��%b�����]
~lm�P"O�T���G�V����j�[ `�""OH�7+Ξ	lH�#��7?V�f"O��r���&�Zt�
�w)|A�"Otr�!V7ɔ�S�'^�A�y�3"OZ��I'p}��g�LG� 0"O�-+�(�.g�*�@���<>:���"O�����W����se
����`"O�E����o��ɇ)��Z#"O<uB&/ sܕ��(N��dU B"Oֱ�#�)���a��(rڑq2�>��j�P"���?}9GH�#p'�0��d�� *D�0���Y&!&��d�ЫF�n!�oWc�G�d5�T/7�3�45V��a�$�(p�,�p-�2}Z6���B�M��a���=st����7��udW�>�xPD��0;
^��$��m�� CɋE����eEV ?�����I���)��2�{M|��
׵OA>��rCP$�}���t�<�E�Y�5��H'�LR�����Z���� _v�ؤ!�aĈ?��E�*��]�i�j7-E0L%~��5�Y��zgC��ks!��;:��b�3D�P�Jg �d�c���-QT䨅�q
��gF�=��*H>��w88`�.�)WܮU�!Й�4`���'��p�)n40�)@��:Cc̦H),��į�jGȩBta�)03�x���>Y�HB���?��E ,,vɂ�U�i�tJSlO��Ol���+
�[P8�¥�@�w�z�j%r���P��]��lҌhg�<S��O앺��[�b�jT+ӓ5c�j���	O�������pC�͢0����0D��?PLy *JA�'+��U�aȄ)D�F�g�`�Q�ϻb��i(�!���y��F�Z�`�نdK�L᥈�? ��v���L��,�.� ��WD�W+��qA�>�O��N�RD޿_��ɉ�$�CN� �$|Op���ȁh�N<����3J�>]�BM�]v}�!�AnV��NS'(&̜1�%7}2I]g��?��f.V��aeLÓs4ajQ�
B�',�Li`��+_���C
����O7P�ʧ��q6^�q)�'PJ�@��'�h��QJ��O�4����g�&��򤅏*-�@�i�q.x�+�)MP���b@�6�D�)���@
5�Li#g B�e�$H-��@ "��A#�>�z��t&=D�HZ��RBr�9d�w�$sՀ9�H&��-A�
�3KN�,�bj��X��I3V�i{DPD���H�@��Ç�FT�R%�zF��+歗�t��Z�#�;s }D�_�a�~�X���l?� H�����>�'��ٲ�.L�M�v����-y²9��'
��PM��X��lh�AK��2)��/߰�ȅ�IFX� ��/���l����%ݚa�&�;<O�x�Wh�#הuخO��'l����O#a��"O^Ac�A 2^(�����\��ɳ��|�nƭY�����H�t�OȦ���a�h�KĝG�ͳ�'W�u����E)��9�ꉋa"Y������'�4X����>YшW 2�yx��4��F��}h<f�AX�ہ���xe�ͺ:e�Q�a��ռ��d��u0�`����`���=P�y��^��n��V�^}}bH�>��JBhR�u�R�r���y��t!�A8$'�s1�����'0� �j�i[�?� (iQ��
0΄C�hB�5��9�w"O���"o�):���/"�n�8F���/�qOV3��Y��겁�p3^pP�ťrQ����/��'rdA�V��>�5ҫnt���G��
�r�YRdHH<�Ԋ\%1;D��G`;KP �dL�J��A:�Ä�p?WD��-bhm�@ݼ>HPq� f8����؃v��4Qe����3c��.�u2g�J�o"��� 4D�|[c��$��b��2xl]�&C!}��zo���B�B�g�Ъ2]?�y��5m�ʡ����<�#3D���!cñM�،���k�t�Z�ǒ�72�'����%&�'0f������y'�wh�� Q�n�T�XV���Px��I:h`����8�V�����*}��`1G*x)r��O$�9���W�X�R���� !���*�قC��0��
5��x� �c
<�B�@d~��0s�r���Y$l6���4 �.>`��m��U��9(����?֊�BĥS'' ��O���ʥKFrK<K�H��(�'4>p��m������N�@;���'A��@	�9yԉ�Ҏ=^�$�t��
���$y��	�iI��H9�`��Lr�����e�>������ ���u�1$�������Bh� ��'�:m��_�f!�`d����	?t�V0�����gy��Ԓ(e,K�lM;i���1#���<A�,�;k�ObcD�i�X���9$�`�R*�0D��0�� Za|� � ��2T"�Y�����Q'�p=�!�ė)m�[��5  ��ĉ�~LeYnފV��`����x�CC9�J,�*B�
���CgO���'��I��N?��� W�	q��LSE��ɜ��#*� l�&��"O��� "Ļ�d���6j�D媒�ެ'H�ː��
s�6u���iTV#}�'8�iZBS�L��3
P*���Z�'~�%����"y�lL�s��QP	�ڢ:�5��*F</l������0<qR
��M&lI6gTU��`���r���95E�,2̀�ҌH*Z��a���4b �!�Nʊ	��8P��I�!�Dڍ6��Ȗ�_*xǫ!��"ZXz���ܮG����e����EJ�'1Mx���)�����1[�Ytv݅�pb1X�D�J�
�r��F3@�$Rw� �T(�A.@:l(+d��c��Z�z�@�O�-��a�>[Q�JU��v����'b��yƌO�`kTq@��Ͻ9����4+QD�0Ɔ����W#�)��d�rŔO����B��<t�W
ܖ˘�hă&�_� t���x��MI̘�C4d���+B�0m�PCd�H�7O|˖ ��Z"��(�(��Ķ8΀�`+�1��$b��$�F�]}(��Ať��� ⛃b�@�������#��}%��`�h���^�yڎ����p"��gL���1mKd\�����&`,QYFdYܮ�yN?Q��̈r�7�Z5�֣gP^������*���	�x �#�%x���
2sO�|�J��6:t����(;�Ej�̒�h���d��4��5
~LD}��N-��A��L��LA�OTh4I5ЌI��heP��QZ�'�p �#!C
_P�#�O�[\��'V��'ܠ{z���Z��}��$Q2��à � 3g�� E K^�<�UAV[rI����7߼��@���Izk�m3Q�����g�6B&ҲC�&RP`��,st=����7@"ҁꝃ���G�����+���=��v%���񄕂}�Јç�@ ��8�ȓF%��Q6��	P���{��_�ObZ%�ȓ.O���Թp���k3b�����ȓ.	����&�� Q3
s�=��r8jq�B��<5<j�(��C0;ⶵ��% 4��f,��#	'DȈl�0�ȓ�q�@�A�S�$�;2X@��?��|���X C��ن(�bl�|�ȓV0��
�ܭP�ְq��_"��ȓ[b��,�D� )�cK�k�܆ȓ	pX�`GNߐ� �(�j۸ن��	�F��`f��l�o�L�h
�'�B�A )V-����b��i��!�'�Lt���F����@f�m��'`P�0@S��6E�t�݀].�!�
��� ����eҷ*	P�"��^�P͐�"ORq82L�<F�Hx���U���z�"ON隂lR:3�ic�P�3�t�@"O�a�ě�,��pp��@�kz��%"O��{���B�\21f4x�1[�"O�e��BʎzB�R��Ǟd����`"OZ�*�RӚ�h��?9ݪ���"OP����
ZBr|CK".�@���"OFA���R|��)�]�k��m�"O杈Ҭ�DAvp�3`E�s�\9)"O��j���y�މA�*I�X��p"O����}��s��8�p\��"O�(r�H��Mb�j�![� �"O�xO4{�.����"���@
�'<��������U�:y��j�'bC��}�<�s�45�T]b�'j@A`]::G���3bڑ ;^4��'�q�UD��g��xC燡l�R
�'�dq�S��9l��W����	�'-��(���#(�
	(�eG/V����'�t�k㌔.�9æ�$V����'�Xl��܂q��U����C�����EWf�:6�%M��H@$��<��0x�-ؠ� ��ȓ2�b�17,��s$`�B���5�Ќ��q����{d�i�y��4�ȓ*�*	9W	׺z$x�&�	M�n,��C�D F�O�P��m���
��P��d�l�j0��92��BJ^<W2P��x8��&�ЫP���Z���f�B;|�'D��Ă(Tt�S�O� �:��C����K [�0�Ҁ���a�f�b> J?c �eF����ߩz�pD�V�1���qf��M����Oq�����T��D8�e��i�`\��
}
3b#�����+�n3�%���k��F�8�M�5r.�{��@~2��=o�L�çy�A�$�5Y����jˇ"�*D�'�Z	�G ՗A�E��'p|��s�Қ��#�a�*H=t4�E� �	�: ��槈��� �ɐk�|�2��Y�+8���,&���HG/!��)�ZA�P	��4Ӫx!�@Ҟ�cv(��hjs-�<Y��`>����e����YF������Ym��TQ+����S�'|I�k��Z �p��C57�|��'�7�\�����ц_j��i�V�?��O�l���]�|�t��b.P 6J܀N֝lZ������M+�FC�t�S*L|�UG�
T[�Y�W�]�:k�u�Zq��`��yӂ���0�ư(�$��JФ��}rBQ��'�]���
v���Ib��'��8yj���O\�b��ɇ��BD�Y>���$n҄!�7-Q�R�@ �G�T��]�������S�O�`�r"E�{ڀ� C7)@"�c6D��1�%(X��pq�;e�`L@�4D��"/��z�H�	!?E�4�Z�?D�<:��=b���`�3�*�)�c)D�X"��    ��   �  4  u  %  ?)  ^4  �?  �J  �U  �`  l  �w  ��  �  W�  �  ��  ��  ʴ  �  V�  ��  ��  [�  ��  r�  ��  k�  �  h�  � � 7 � � M" �( <2 �; "B aK �T �Y  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9��CZ���1.*��5���#D�������=9js����]>+-B�I�L,����ơT� *S"0G��B�I�<w<̉@���R��Xrȕ(Uv�B�	�n�t�hՈ7Cn���ӳ;�B�	x�Ψ3�E�V�B�ʑ�ޕ-bB�	�K��� L0B��h�'��O�`B�I~����b��L�5��£~�B�	�0�dq�  -Nz����� 9�0C�0>a1%
�y�N���.M7@B剖+($�w������Ο&|`!򤂰V�dS�D�
��PZv�I!��"���㰁L5=�����	�!�ӄA��a Q�&�ʀp`�0#&!�$\(�����N*�Z1�f��+%!�D�J�ݨ�H�UwP5hd�	!�$C0�d��#��1a��ɷ*���!�$J�gÔ�[��,;�2	:D��J�!�d�c�\���HOOj��q��o�!�R 5rZ@
T�� ]VH�RbY��!�dI�{g)#��MF�EQ�J�7_%!��= G4i�� �<+������5�!�D
�[�T��"D�*��Mr�N�2w!�$�aFڈ�&�ذM�t�D��l�!��.a��To��6�F|��,	�v�!�DQk�m�D"��W���wN@h�!�X��1R�/߽`v�S!/Ìk!���/uӦ&�(__�Ո!�ǖE1tܙ�I�X�Ļ��̓�!�ԉT���k�E[*E������6#�!�d�zr��h!ꖰg;l\��cT�t!���k~�X oF>@����c�#�!�8H�Lk��7�Fxk��R/�!��Z�^l2��^ a���Rf�L�,�!�$�� .!���"S$�*�.��2�!��0BYڨp� �:8P���KȝW�!�*@�X�Oފ?g��ॠ_�)�!�$�P��+D����z�� E�!��  �!�O�M ��#Y��"�8#"O<��"��5Jf<a�AmJ-�Xt	U"O0�8��+��k�삓���"O����HM6��JB1[��ЫD"O \�!�Ðq����g)B�6 �@J2"O��FG�`:�}�C�F#f,�3"O
��'ME:,�qq��s�(Eg"O���	�;y�t:�ɂ��)"Ov� 7�	+N�H ���K��� "O��c�F�T�ʁ�Ҽ'�Rx�"O�t�䃋1��xI���VfRYj�"O��KU�_�(>���!މ�t�b"Of���m�3��P�N(8���a"O�J�K;kм�2R�I�Uh�@#"O����_�QbKZ 2�pq�"�-�y"#������O�sd	���J�<�SN��M�غ&Q���9Í�y�<�Ed�GW
�f�[A'V�vd�\�<�㧗�E�����8��3&U�<��M�*%(0(�Vː�@3��Ӥ�v�<A�C�{c2(HW���>I(�)v�<I�_p� �S7�эF$�4�4m�t�<�6�Ì�8 �%�{�$@Fiu�<����6D� ���υM)	��p�<YOB<u�N�yt�@&t��(0��T�<ag'\�*�%�fW�:�Y�fmEl�<1��2�(a��N�9�"}`�
�p�<����Z����(�^�m�S��G�<-����bA�E�� ���_o�:B�	H�΅���b��y &�*|B�Ig��X#�'cz�`DO؛t?B��1V{����ʑ*O$� *(�B��#)b΅1���:X�Q�/P�3NC�@�j1r�ԈS&�mSG�=X�C�I x$�A9�2?\����όv�B�I�o����7�ю Kt��GB��"aC䉇+J�;���:~$ *�C��S��B�	��0�3vӤ2�*!� �)��B�ɫx8�l�tB����Ԛ��p�B�	�VV�IP�MK�?�@rFY.!�B��;2?��rq��:��4�6!ҵh��B�	�s��*�F�30z���/Q2k�B�I�M�l�8��	)���q�[�B�ɽy�Zp�L�	p_�4y�$��]@B�	�B��
������r)]�~R�C�I�O�FT��K����RU�Z�͚C�I0#̓ �¥ 
P�qW�T�G��B�	�M��{�E �jlDp9u�ǵ��B�I�CJ��Q%�Գ�bH:ņ@�?JB�	.?_$���ǉ@�~%:��Ql� B��PY)�r�A� "���iܽa�C䉻>�iQ�-�Y��b2�[Y?&B�	�9���ʄ'6"�����	B剓KhZDJ�"�+H���$�F�FO!��v[\9 �&Q��t��$�̺H!��9b�+������$��
5!򤘊bE:@yb�+��r%�U5!�dX3m��t��^#�̤[��O�!�$��\�J͐�J́*~�{�$F8,�!��$�0'����(0�ڻP�!�dȠ�H�ʋ��(��
�!�	*��4A؊k�$�"Y�^"!��Ime�!���\j�r<�5�Y�<�!�$;MM湈@W�1ʦ��nI�G�!�� p��ˉ�	>R��t�	,J�p�B"O�9IU \�`6� ���Э��"O��kNk]�9���97��8PU"O�E@f$��bk���fF��t��8�"O2T�.� ������Ρ7���YU�'t��'���'��'���'���'zİ�r)�7B�*�����) ��'�2�'b��'>��'���'�2�'��R�i�F���*��ġK�T:0�'��'G��'��'���'���'��QJc�L���:C�T�OB��s�'9��'o��'p��'"�'E��'7��0%i��:t<� ���J��y��'���'���'{��'��'b�'�U��Ƅ[hj��d�,"�u@C�'pR�'���'CR�'~�'��'~���G+�()�a�5���,(n�X�'�B�'��'f��'R�'"��'�v�R�Q0A>�k�U>OA~��'�2�'*B�'���'(r�'K"�'�lu(����[i¥�TB�)������'wB�'���'�"�'�2�'��'y��AR˃(@�����_�}5 ���'���'��'���'�r�'?��'�@���HJ�V�f����O�]0(�'�'�"�'�R�'�r�'���':��'���w�Q����&Q�-7hT�P�'H��'q"�'B��'���'=��'F�i�Dێ
_$x���ַ��Uy��'k"�'���'+��'�2�vӔ���OR�9^��		��=:~V���[y2�'��)�3?y�i �MBŨL<u���Y�I��'��	�T�?�.O��d�Z�������+-���)���i���$�O�ph�h�J����j�H�Osxk�&��qB����훸:ad=C�y��'`��Z�Oz�8���G�z:�偰[;<���#�>Y/OV��.�ȟ�]�K�`�y�i�6�^���d��?*�E��ϟ<ϓ����x7My�x��ѲY�vp����(�X<[`�j��J����s�����'"�Y"��z`8� (Y��Þ'#�I`�I���O"�(A�0B���P+��ĤD�,�O�ʓ�?I��yrR���NE B����`,�j	е�B�+?��o�f �ťT�'o�d���?A�lY9_�t�*#�#��!�����<)�S��ycE���\�J!��œ�5�4U	�_G�Iy��'��O�[XS�H��4`0��C��
`G�$�O.���O�q2V�yӺ���4!��bMQ��VF�!���Dd؊fL[��䓀���dZ�@��IA��!9{yY��]�I��D�O��$�OZ�?��$��\�D�e��f8/Y�%a�	7�M�%�i�O1�lX�AlO-�$\IRF�&��AIb�w6��*1�<1eV�=��İ�䓆�H�:1�m�wf�=W3�,�s��#&a|B`�>9��prFcT�s��iP�F�9A������?)�"\�(H�4Q
��!|�NM�O��~O|]����*�;S�A4a��6-h�p��3`�*�P�O��Ж'��4�w�D�R�.(C�X%;'f�a2���'���Ud��(����*^�}��C�r�'��͸>�O�ҝ|"��|�P|�4��;nи��)G�jO6�lZ��M�'� h�ܴ����	�~t�`� C,8�!`H�.��R����?!0�#�$�<�����+gKʟuc,}�`�O���'�B�'orP>����@�s����|H@�[�%8?	/O���O��IU�'h�� 1욁d"������ mN�P�F��	8ى޴]�i>8��O��O��p�̍t���;��`��X�Od8nZ�f7b��vj�0z��@�x��Iʟ�	ğ��?Y(O�0oڰHvJ���ʍ�}�QjT,CJ��ܴ\����$Nƛ֚���T����j�nyOA��$a���>F���A�e�y"\��	џ�������	�p�OLDp�V�"'�j���!A�JP��@�>��?���䧮?�Ӽ3�*��z�`1� ��y�gS��i!��O��O��E1��f3Oʔ!׆3�\��e�W@��2O��5���?Y�(��<1���?A�陛*�2Y���_�]�>I	��؂�?Y��?)���$�a}r�'��'�bA���;X���k��K�4����$�<Iֱi�7-WB�62=��ACL��,��9 Em�*3��	֟<ɲBY�'��2C�ty��Oט��I�G�r/�?)unѨPN�`����՘h�2�'���'.���X� T�p\���ʝE��U�q����lK�O����O���:�i�Q�T�'�D�ڑ凣A��Rv��y�4}:���g�r� Si���D?���������3	�F��T͋κ���6~��O`ʓ�?���?����?����Uqv�		�:I�T�ݪ.��Y(O���'^r�'���d�'c�"�jZ�W�D[�E�Jm�`�W�0�	ȟ�%�b>	KT��7m��D_�NH���L w�	spF>?��#�F!����<����D��lB~��E�B'	A���o��G����O��O��4���5�I���s�V�!�l�4�F@���g���In����$�O��$�O~Ȇ��B��rB	P㚥p��A��7�6?a�B��	$�S��� ��jcI��m���2��݆Kg,,�g3O��D�O��D�O����O��?�s`��)h����G^=~z��C������ß���O��O2��6��0;f�� EJ�Lx�����## �O���O�� �Bm�6�.?� ��M��x���#h�>���V�@���d��On9�N>�,O���OV�$�O�t�p�ȓq�^�CP��9��͑ĉ�O&�Ġ<�S�@�	�� ��y�d�|z���A�Pĉ��d�����<Y��?�K>ͧ�?q5E���IIREV�sB�CiG�tS�:
Q�4Up�'���,��:d�|�N��}�J<���6����K�"��'��'����[��ܴ_;�����LV����K���$̓�?���?��T�|���ڌ�G�%�%�����p���� �&�����?Q��2 B�)RO~�'A�C0��iD.�HQ',�yT���Ο���ß�����O�xd����_,RX ��y�@��>y���?�����<!�Ӽ+��O�k#���txc!+���?������|���?��49l�<I4��/�LxH@�Ȑ>��m˦���<�H�U��d�6����4���D-0$0�cFN�1���k�-,|�D�O����O<� ���p��̟T�!S�I���5$0����Pd����O��9��Nw�~UP���")�\� 	�/����?pR��G� T>c>݊��'^>��	�Z�ኤw�$ەH
>�D8���' ��'���'X�>��	.[=��U	�(��["M(<����	���d�<�����yg��1`�U��G�=��ܻ�
���y�{�Dlo�&�M%��Mc�'R�L�+���S1.��ʵ-KO��Y��I3'.b��s�|�S���	�����؟d�IߟlpI	��=�jK�B��ȈJy�Ȧ>q���?����'�?�0�J�|C.	q��\.0#��c@����OD�� ��O<��O;�-��CU�7��-��"܇bV���]�T��[�`X� v�"�l��ay2��1έ�PkҧY�𸓂X�Z�'���'��O/�	*����ON� VKKNAu�!,M�k��r��O��$0�ITy��z�Ƽ�	Ȧa��e´A��I����i��X��#����o�[~B�C�<�lL�S�0u�O�g�I{J� Q� �fH1��Գ�y��'-�'���'c���R�w���Gxf�8���Z!eW&�d�Of�$�q}�Ox2�':�'��I�4��fjnŀ��H�5�
���-=���O��O�Qմi>��7t�.}hg�y�={�+u����w��j�q�IEyr�'O��'2�.�<LЄq�5���q�~p鱣ɕq�r�'6�I���d�On���Ob�'*E8��W�z���X�&_�NB�`�'��Iߟ����S�t&F�JE�"uҠ��zAWReb̫�J,P %Z�[���*�2hEm�	��৪�p b�	�i�	ȟh��ӟ$�)�[y"Go�,)S���XX��	-bMļH�6OF��?�RT��A޴P�.aX n1�Hp;���P��
��'��F��W.����< ��Xj+���jyR����[��/en�$��h]:�y"P������Iɟh�	ҟ��Oޒ�*�M?M�L0�������)�>����?����'�?9�Ӽ{�I��
��l �b,A8��ʦ��V�ORO1����#iu�*�	�X�1�W;�,y
���7�@�?Yx٩C�'C�Y'�̕'��'&`�1�#�d���Hl�^�2t�'{��'��Y��@�OD��O�d>Bq���.Q8��70t�㟌�'�:6�B� &�X�Ď�$O�x!�-�:DQA3?�Bh]�J�v���%��N�b����?q�9�^�U¤j�R�åE!�?9���?��?َ���O-�JW5Nk][AHT.{�f�S��O�u�'�"�'���4�`�ˣg]9ZXڂA�
���1OV���O���Qo?87�.?�f8hŲ�i��	c� �h)���$шb�D�H>	)O���OP��O��D�O�5 � 6���&R�ח���m}�'���'��y��#8�Dp�C�È20lb �շw��	��@�	F�)�>����=Hf�؅��+�4lY�Y!�|�V�w�{��f��O�ʓ�F�C��N=l�J(�(D������?i���?!��|�/O!�'&���B���F���j�^�թ����'"�O�˓�?����?�a��s����:F���M8H+v�4�y��'��7#��?M#�Of����% ��O$-*����� �C>O����O��d�Or���OZ�?]�!-�@�(��TL�4g�M
���ğ��	ȟ� �O��͟�$����.Ó{v�%��1��u:Ԩ	X�	�t�i>�XPaʦ��'c��0��6b_��c2�M�<S���f#�J�Xy�����d�O��$�O���O�:������	�#] 	�%ڿx����O��I���ڟ��	�P�Orp٣'L����2��;[TdX�O˓�?����S��EOH�{'.Cs�r�˂�U-v]āAq�1uқ�n�<ͧX���l�k�"�HsC �te�i��Iuр(�� ��ڟ��)�STy�s�86վV$n
����&q�<���?����?9��T�p�I�`#h����7`1�=��G&t�	�|�N���a�'�&��1-X�?餟� ��	c���v�l8�] #5��S5O��?����?A���?I�����ɹglД(�h�kpF%@�/°/O��'�r�'"��d�'
�wv���,��dKr��#im���ia�'m2�|�O���'�|%�i#�V�}lj
1�#7���*�Fܙk?�֡
�<8R��7iƓO>��|
��vdjE/?6یȩE.V�a�I��?���?�/O���'���'r,�6����+�BAzn����O�˓�?����ᖽ�I���'{8&\r��@~�"��O���Xֵi^��~5��'&�ؓ�(QeH�M��}i� @�ko��'���'"�Sߟ���
�6�z�����/�<�	��Zݟt �Ot���O��$#�i�����߬��E��(��v�s�Ds���Iϟ�̓1<4mZ�<���>����j�?���I&����j#x�����s�Icy��'���'��'��H��X����Dj\|�S(�1_�	����O��d�O"�����E0,nݐ�G��h�%�/",j��?����ŞFTz�p����
:�H�ẻ+��9
�����M��Q���$��=���"���<��C�l<Zt�5�Z�
Q�WD?�?)��?����?�'��Vt}��'�P�c�]H��ّ���&�P�П'q"�D�<Y��?!����I�.Ҳ$��|�1����Č�����M+�Ol\�2N��ڌ���w�b���(�8B���b=!����'�2�'hR�'�"\�b>���S6��Qf숌Gi���w�����Iݟ�9�O�	�O��.����5V��X' <@<$u���X.c��Od���O��1l6M&?q��%�-Ɋ��0���ڎm ���O��`I>)*O�i�OF���O����D]+bX]�S'�>c� |�t��Or��<rQ����矨��@�4ju�Ì�7�ع��	�Lt�'u�I��͓��S�t��1Dw|	�,
-3�.=S����z��CdK�X���Bs]��S�xB�w�	-(�9�'k��� 37nԒ?���Iϟh�����)��fybc�Ё�F��$*Np���DܲC�-�t?O��d�O���1�Izy��'��"jZ	:xy�A L�T,��	�7O�7��uz6�4?%�����iG*���_���-p`V/,��HK���<����?	���?i��?!*��X�Q'��)Oȩ`ч�Sx���G}b�'�"�'~���4�80Q�:`oh����˷$�T�9P�KӦK�4[����O�\y9�i��ėARX̹bOC�iq���'k� �Ŝf�
��x�`�Oʓ�?���U �%KU �<N�Q�QM�H�,<���?A��?-O@5�'u"�'�b�U"��l����sd��1VjY#s1�O|˓�?����|�hh՚M L����:!� Y��?��\�{����4l�I�?�[t�O�d[mW�Q�ai�y�(���␅S"��Or���O��$=�'�?e�L<i	D�c�'B6��$:#���?�T���Iٟ��	d�Ӽ#ЈƕtJ�9d�Q�;�����<I���?���RO���ٴ�����B���F����ND�sC�f覀�t%�����d�O����O�d�O���Z��D�[��͘���z� ��PQ��+�Iş�Iʟ�%?�	;g���kV[~\�I��
%>��ܗ']h7M�ڟ�%�b>y�2���cyPy���}��Y�膈Q���:fǔuybfE�8L�IS��';�Ƀ6�B��FPu·$�FÈ�I����	����i>!�'�`듅?s� S�����ٌ;m����Cҫ�?����'��ɍ�M���'���b�%y�"�_?.�i��SS�d�s�i��D�O�xJgꆉ�rD*�<�����ӅT*#�|�P�TpULt�r(Γ�?y��?����?���O�^��!� +�Hϔ^qN��p�'���'�d��|B���?YN>�恋#V���SW�t����a�l�'��z&�Р�M��O�y0��B	5J�m3��O:$�!c�Nt�>� ��O8ʓ�?9���?I��p����,T$"�^�������q��?i+O���'2��'�BP>qs�+��Q�;�oݸ!�}8��-?�.O�o/�?	M<�OH��ƒ)S�LLg��	7��epv��.p����vN�i>!��'S�%��[�lQ�d�8��B$X�y$�Dꇢ��T��˟��I�b>q�'�7Z�.͒Ÿ�a��h��l��B�u���Ot���Ov⟰�'�7���R�@e
���z���ĠWE�m��M[�-�;�M�'�BjS�U�d��S&��I�I��,�W��e��s��^6X�(�Ry��'���'S�'��^>�B�� �N�a�G�;�Ɖ�3����d�OF���O��N�$�O��F=]+ ���	]� Yѭ�%yM���Oj�O��O2��B�d��7mh�0ZAl��z���#G	�qm�1`c%d�L��Jݸr��� �D�<!��?��E�Q�XX�-N�0�pv�X�?���?�����D�h}��'��'	*0�S��LWl\(� �x֠QZ����<����?YH>��Ǌ2:TıVNŢm����ǯ��<Y��M��,���6�MeU�h�Ӂ5l���O� ��Η3������ �z��O���Ox�$�O��}2��)��z��B�u>�89rkM�E�)�b���П ��̟4�?ͻ`���DK#i*x� t���.3"L̓�?���?1�ڟ�M��Oݡ�&����� :|�1bPr��u���'$ �mK�"�ģ<���?!���?���?Q��^�5>��Y��r�&@���$Pl}��'��'���y�Y�c36 `�bW�~ �hS��]�E��	3�M��'퉧�O�L= E`�!�ɀۧo�e���L�7A�!bpQ�$p%�	0Vr��G�Iy⃕�Cb4!2O#h�֠A�U�2*��'�b�'��Os�	���d�Of��Ě�0�,�s7��:�dP%��O��$2��vy�'
R�'��X˳�;`�X�B�-`�� �-ՙ(���7O��E7�2A��Oh�I�?1�]p����!lY�{����Ҫ^�.�	ߟ������ܟ���`��DR��V9f@a��[�����?�4$�i>������%��o[M�h��&ȃ�h��I`��ӟ,�	������=��?T-ֶ1H6u�񢆕�ࠈ� x�`Ͳ�䳟P$�ܕ'B�'�"�'J�(YƭA��D5S F�$D���'�b_��Q�O���O��d�|���61#jAQU�� ~��P(b~[�d�����%��'�1�I�#M�6%�Fm��Z	����7x��޴C��i>ᑀ�O��O��k6CT�L��2ti�)�Պ��O.�D�Of�$�O1�ʓ���f 5`8��j3n<nulES�Ȅ��y�S���	c���$`��#5o	�Txb���X�I�|9Q������nzK8�9n�p~��V<�h��'f���>N��P��ā,b�0ف�.V1����Uyr�'���'
B�'*2_>R��W)s� �KR��$q���!�0����O����O ������O�H-��Z�dݩh����\
n'��mڄ�?)M<�'�*��!v5hݴ�y��]	>����C9^Z�4���yn Qr4���0!��'s�I�d�ITi�i�Fj�х�r4����F�˟���̟���Zy�n�>-�Ms���?Q&@��ƈ�T'ѩ]5��+�/����'���ןX�In�5�֭Ц`؊t������G�.���9jp'���M� ����Nq?�����X �&(��Qe,H7_`��S���?���?����h��D^�J|Y�%���w�V�1��N�
���$�G}��'u��'��O�.=rrg��+_�p�H���z�$�O��$RΦ��Næ�͓�?ѕc�R|��ɝT詪g�J�.��pp�-6���M>)(O@�d�O��d�O����O�!S���;Q��f�W u�>ܣ.�<��\�l�������t��� ʱ�c&��Q��7	*t!�fyr�'?�0��iE!?{E��'K�����3w��)w�X�K�˓�h�����O:y�O>�.O,]�����+�I"���e�����O4��O����O�	�<yAR�H�	6[%d��Pe�8)֘zW!	H_b��ܟ��?A+O�o��?��4=Ҵh����#r�<��" _�^¶9��{�ٴ�y��'���9'�?�y�^�,����Yh�B8Ǭ�4�ύEś��g����ڟ@�	����I���K�q�]�4)[�w������K�?)��?A5X����(�Ik�	6
w�xruK͒\��,bV�	O8`�H<Yּi$"6���3Ă`���	h��DL�iԪt��
�1\߼�{Ql\�8&����'�p8'���'�2�'�"�'�0U:�ӁSP>%2��l7�����'z�P��٬O�ʓ�?�)���:�[�f�b�A���WfB(PG����'�6m��q{O<�OL�	`E3+�B�@�&(��HÅD��x���+�ca�i>%��h�;cj�'�ٲq�E&t��4��Ӟ!����' b�'d2���OS�I-�MQ&Уa��Xg�\�k� ��e���<.O���6��vy2�'��@��E�4"�zqgዐ�Y��'jb�T�pG��0O��䊘sD^���'$���fQb�ʒ%W+\0H�I���gB���ly�'��'���'o�S>�:�d­gz���l�kU|�[`k�����O����Ov����O�N����t�Ⱥ�Ђf��X2����O��O1����r�x�I�Xְe��e3h �]�p�,�^�	�Yn��F�'�P�%�����'�|��� @�d�āhU$���"���'��']"Z�TA�O��d�OJ��	�:]�u���N��'��0�⟘�'�R�'��'��t��Ɲ�6��R��)q�	Ø'A�Q�,_�A� �2���?Y��'�,��ɣ.{��b�b΍qqb�c !�;q&L�I⟬����8��i�O���Z����������,��0@�����>���?�����yW瀸G���2��׀�$@`�ֱ�y�$l���	Ħ�;'o@Ȧ�'� `�@�?�{�i��ª�1�-ˠr���)M ��'�	�T�I�8������V�����k��I�Ь�����'Q���?a���?�H~z�tZ�9�˚(J����K�Z��*�O����O�O�O��s��+	\^T�a-	�W� X��M��<)@��@U���"��t��CW��ty¦	VD �BG����T�K:r�'<b�'9�O�	=���O��Î]&U�qACD�Bu��>O��0��yy��n��q�	�12����*�$ �%�6ݐ@.܌y�6�n�F~RC��p����ӣ
��O�w��k荫BIz�ٓ����y��'�b�'s�'v2��9�8ڴ�'\�X�P��_���d�O��D�]}ʟ���=��Z�}�"��B
�+�:xфE�֨�$�|�	Ο��E8w
6�=?�#Xu�? �p��ӴT�.ȇ͗5V��r�̊�?��3���<���?i���?)�$ĿUJ<���C�3(\,i�Y-�?�����a}r�'[r�'L��<�1����&�дg��v�`����������S�����6�����;3`� ʴA�h�(h���*�`�C�V��ө:��MX�I$v�Z�G�X�b;�댙q�A�I�d�	�p�)��dyr `�T��0��c%��c���zI����5O���?ɋ�X�(s�4[t�0�EJ�<&�&0���V�<Ųb�'��V�A�E�6���2�G^�x���NyR�M)n$�M�"&�zI��fR(�yR�@��˟��ٟP��՟|�O9��`G%՜i>h` e�z��9��>����?�����'�?	�Ӽ�� ����+S���j�����Ku��\$�b>��)Hɦ�̓d�U#����KF�k>���pd� �g�؋F���o��Jy��'��Ŋ�*F�3�ٍ]�*�[׎ Sn�'���'�剐����O��D�O�P���˔z=��0�^#F�^���-�	m~"�'��V�1�D�Nv`�Xv�d��w�9V�x�J�O���!/�X�L��u<�i^��?�ub�O���jA�B�n�J���,B��iJ��O���O���O��}�;E<1p���)㘀� %���\ 0�Ga��ş��I�0�?�;`'H���a��D�p�ׇG7~���?y�4��F
?�M��O8T*�!�
��X�����(��z��IȒO�˓�?����?���?���EsΥ����9elR��[�F&P�P-Ob��'������V������ �P��=�Ă[*����O���2��)H�jh��R�ª4�b쐆'J�E{�Iu�V|�'P�,�a�j?�H>�(O`Q�(�}^	(���:�M��g�O����O*�$�O�<�BS�����XΜ��#�ti�ٳ�m_����	����?9/Ol�$�O��Ą�4���H�
ʤa̒P�FD1Ѯ��g�p�@�DD�q��?a%?��� ZG��ڕh�'�r���	!<]���4�	ԟX��ȟ���o��}�s&�ÊP���
T�S~+��b���?i��g��i>-���'�t0$f����Aٵ�n�%RN�G�	ʟ��i>�1���æI�'��!�,B��ѓ��
r'�`u�^�1��"��'p�'�Oq��'l��' �];�J*i8e�e��U �,���'lR�'A�dӖ���OD�$�O��'��XnO�i0� ]!�"�3�'��6m�O�䟄mZ���)�|���v��(!ş�iG�����1K�Xe�"�tȚud�-����  ��&���OZ��d�
�+D>� D �`T��O�O���O����O1��˓7 ����v���s�� �l��x�ƥ�y�[���Ie����$�ǦyZ#��3����v G�W�<C/�?�?1۴޺���4��ĖU�@qk�'i�˓�������\BuP��ʍQ�"����d�Oj���O����Oz���|���P�X�
#D�A&� �5�H:"��؟����$?�I���J� %�P��&����m��uj�a�ܴ���!�4��������hӘ�Ij�!��
�oV����	������'�fI'�ؔ'���'ĺ�م�� �V�Q�BL� 3��'J�'�^� ��O0��?d��Q�NX�uO�=üJw����'��8�M�g�iy�OJj2�V�5IȜ��1�����S� ���LbD/�k�8�/�|�"�F�7:�L����h��Jן �I����	��D���'3Lx ���R���+�H�F1��'����?���?��w��"��62���F	j�hd�'��7�D���A޴O��q��4���2_�����'VBq�$�	�4� i�s/ݫj@���0���<)��?���?A��?�0)dΐ����A�S3b��k҅��$�]}�'1B�'��O0��5Q��x�ͮ��ē��D�	��M�i��O1��ly��ʒ�/��D-�̡W�L*Q����7 �n��I�33D�2��'i��'���'4�:1FܿY7�#��P�I	��jv�'�'����S�xk�O���)��2�I�x:=2�L#K�����O<�\�'�r�yW�R=.̈�臆� Iݰ��V���S��Ӣ�i��	F�Nţߟ�������b�̛&���2�uz&Y'��$�O��d�O8�D�O��D$�Ӝ (ܑx`i	�H������;q@"��Iȟ�	*��4�F�d�OD�Ox�`c�U�BIsӍ��E-6�[!(!���O��4�i��xӦ�ޢ�0�fJ'Aܜ���l��+?̵:�;o���W�\y��'x��']" ݻ$?�)�dl�T��h���߅N�'��	6��D�O��D�O&�'*�D��1G��N���jl[(���'��Iʟxn���S�T�ݤi�t(�RG�R���?DQ�%�����.�.�	$^��S%S"&Pz�Ʉ&�c@�d\4��T�J��0��O����O����O1��ʓ(�Fo� a�bH3$�0�,�]���'�z����'��	%�M�w�a_R���M��:+l�ǧǘe���kӾpa�c��	��2O�o��4��|y��S��怪&dL�H�>X�����y�]�P��������`���Oi�5��ge�r��>�By{�b�>9���?����'�?��Ӽ��Ƃ|�0�.��\����bj��n��M}ӈ�'�b>-c�kBϦ��S�? d8JbKI�IA����ힰFrnա5O�TJ߬�?A$�7�d�<����?���߫`�t������W2T1���?1��?A���}��'���'�����Z<ŸiXD`�?V�� �B��<aD�iE��$'�Öy�-s'(�w�j�F��I�I#xgF�2!"A| �@$?���'�d�	'8U��o�lp��
���+��0�	͟@�Iៜ�I@�O&Ro��1�p=����S�(�j�!��(��	�>����?q�����y�ƕ��Z����H2���%����y��uӖl��M�c-	�M��'��]����2�3��O�9[>�C!*�e�R��s�|rZ�Vjӆ�d�O���O��D^�7��2z��V��Y�*�+]��ЩO��$�O�$.�I�O�U"PDԛ:s4��֊�.Z����Ǹ<���y��x�Oc��O�59BA��$��EgNJ$u�ώ�GM�ʠY��ptN��:�R+�d��~yC�5h�5��cK -L��k0;B�'R�'��OE������O�}j���>ʊ4��F���FF�O>��(�	Ay��c�����٢T��jL|{!�����;��ϕ'���ll~2��8>�.���_��O��#lU�1��o��Mv�9�*��yB�'���'���'2�I��H?���#�&�\�{�h_�.���O
��o}�O�"�'l�'��yTh�4@}�{��C�	 ���3�|��'`�OJ� �&�i��	(;/�-��mx��	D��ACrN�j�~�|rW�������Iӟl*���P�r�H��n��l9�����IZy��>!��?1������A!P���
6�U��������wyBgqӜ�m����S��+��L�J��F�ĺ�T�)��貲�LѤ,�^��S�m\�h�y�	'��2'�u�(:�%��kw���	ȟ(����h�)�ny"�`��CD_^<Fɛ��?nC\��3O��D�O���5��Ry"�xӆ�8��a�0ر�
8�j�8�cɦ�@۴%f�<2ٴ���,�:<����~˓O��ܡ����S���V�<te����O����O���O���|�a��rM�a�/��-�����>.���d����$?a�I��]d�.他hȒ|� ����Z$7��TI���ٴ$����d�O�)Z�v4O�u:Fb��U>=�u���/�,�Ɂ-1b��'�f}$��'��'�����J�v��$8�D�O�p5�'�'�"�'��[���O����O2�䜆3���@�-�6;�&h���^M���'!d6-���l$�hd��6�C����ᇅ(?�O��,SX�Q�O���+PL����?�D��" ��G�YV�xQ�	��?q���?���?���9�8g�A�Z��PѢ�QրP�f�O���'w��'T��4�b�j#JE�$��d���_D��t�O��kӈ l�*0Iok~@	"lVl�Q1J�x�L$X�6��өVP��i��|�Y������ �I�(��ğ��U�PB���e�0A�����h�iyb�>����?���'�?Y⁌�P��	��g\|�35�M��$�O��4�4�����O��{'��F��܊�� kO��Y�_.�7�\y��Ίp�pq�������ԧL����+t$(���B?�����O����O��4�
�B;��蟨�6AՀr��U��A_�~����GF�P�Ig�����O�d�OR��"� Mp�����v>� �!_?�6�!?3 �^En�l����{'�ދ/jfR.�/X�ƅc���I��I��\�I۟����.�G�t݈q��#u���]��?I��?i�T�Ė'*R�|r/`MZ[�痥G��	hG�C{�fO(�o1�?�Ӆ��1lZ`~2/>`8�}e��~y^�;��֛s��hH "ğ��|R���	�T��ğ�:��9F��u��i��]rƝ������P��SyRB�>���?�����iƑ�|��6me�H��J�a��	`yR��&��o�)� �t�t��"��O|nU��F�.�ag�S!L��,O���?I�3�D�+�P��h��*m��OE%?���Op���O���ɸ<���i̬p(^�&o����̢,<]`�'��	���?.OΜm�*z��KQ�]
���N�
^�Y���Mf���M#�O���nD�:�j�<��B�O�.�" ��
a``ړgH�<�,O*�D�O����OF���O�ʧh�N8x�S)K@��8�ϢU&�X��Y�L�Iџ���v�'�?ͻ-�60�Tj�T���@����L$�X����?QM>�|2�I��MÞ'�J�:u�C�����L��Б�'F�p;tjx?iN>)-O��D�O\���@�W�`�r���#:U�R��O��$�O�$�<yY� �I����	� �"�j�'�Z��Z���6>(���?.O>���O�O4@��� ~�T�P(W�?. 9�Ж�h�@�?m�s�a,�Ӈ?ia�Ɵ��r��|*4q��L�M�ޙ�@�Hǟ��Iߟ ��埠E���'�t��çØh��u��L�p�v�:q�';���?���?��w����W�7Y�rXf��~'"}��'�7���ܴH6�Xߴ��� >�rH��'\�H @q-��w��1ɑ&h��K`�%�d�<q��?���?!���?�:V ��5�L<����-V7h�ʓ�I����۟�%?����=jD��dO,K������^�;b�'�.7-�ݟ�%�b>�i-� ��yV�L8U�x�"���ݾ��K�b���/�>t�b��O��3K>�*O��F�I�^��@���z��,J���Ot�$�O`���O�i�<��Q�0��61��Z�E��5���d��>ABd�I�,�?�-O�In���?�4;�f�P���O�ti	�D�`v�� ��M��O�u��ϣ�:��2����P��`��0ѺMS +ۑ2���9O����O����Ob��O��?�9V�ML(f!s�Ӧb����'KRڟl�	�lk�O����d'�Hȁ�A�`m`�Ε/L���;�D�ϟ�}��	��@��64?��hn��z�-�
B=����O�$�+�f��4$��'��'�b�'����g�;�V�1d�ªS�7�'4Z�T�Ob���O��d�|:��_�AT�QT�9rT!�B~2Y����� $��'\#*D+��πf��AA1j��=��5�J4r0$�i�4/ �i>ɋa�OR�O�H8��UZ��SG������O���O0���O1�p�Z��ȉr����ɟ h\�ţ	�y�P����O���d�Oʅ�W�ؚh�0�'dP<p�Ҡ���O����Yo6�=?y������I=��Ǉ?n蜙�Ccؕ��g��y�^���Iٟ��������ߟ��O�ܤSv�H� \��#K�w�ԍQ�ɤ>�,Od��:���OD�4�
��2HW&wz`��fa΢ �tAs�Ȧi����Ş
���kܴ�y�I���4�' I�U�l�r�F�>�y*I!{�8�I*gc�'�؟��Ʉ]Ҹ0� JBf:y�5 �'<k�h��Ɵ ����X�'X�듃?����?����*b=Pl;!�\�(P�9p����'U�		�M;6�'R�'>�b�%B�"`�l�ĭ�~$����O�x�b��+�N���&��O�?���OT)�Zo}�`hW�"<m� ��]�?q���?����?��)�O�0�D�1���Ѵ \>`&����Oʤ�'��'�b�4�l�HӌP�-k�`1W�>�n�9O�]l�?�ڴ#� �ٴ���חz�\��'3�´��曧eo"��n�D�j�a�	-��<I��?	���?)��?	�^�t�J�Ň 4� HX�O׾��d]D}��'02�'��O1�
c���#A�0�x�W��,���M��'Չ��O4�p��� �<\�����)F.`��+x<�sQ�� ��6E��G�Ivy�M��1��La`�^�40fO�f���'���'��O��	����O2�F���<�����,[�X��S�O���2�I~yB.v����	����'
<L��J7���&�������7�0?�w��/pe���R"��'���℈\�+�CT)	l$@����<���?y���?a��?����F�%�D�����F��|�U7[j��'@ˤ>�'�?�����	G�ыt�O70����*N�Q>�ْP�xAu�����`5��|��G��cDާocv(�W�޸U]z���͉ +E������䓪��O����O(�䒫m4�,���\���lw��vj��O�˓g�	Ky�'���/���B%�G`�5���_W����女�����S��ˊ�1p���$��3�d)��ۆ9��X��ʃs���@c\���1) ��s�I�,:,�k�Oԋd�0�D3Mgz��I��d�I�\�)��ny�)b�,`B��>���Ó�@Sf��g;Oʓ�?���X�X��s���ML Nv����C�dEh)�	������ئA�'�D�c#��?E��@R2�TY[�AHB#A
v<��34OH��?����?���?����U�.j�=�v�9~J(�bE�@�ק��4�?9���䧓?��Ӽ#�*��/��a0g��k].������?����S�'}����4�y"��8�iQ��&X�B,��K��y���(�}�I k�'*�i>��	�E�R�zv$A)�� ŤP!<3��	���Işx�'���?����?	
�=��h��K�7�N���Q���'��Ɵd��Y��{�6���H�~�Ƽ�cL=?E��^��1���?~�$�|Z�"�O�$��@>9X�/� #a�,��:���?Y��?q��h�h�d��>�i��A%%�R]����U��DKK}��''�']�O�n�:JUQWLU�Ĵ���G����O��D�O�s6�}�0�5m����)���X8��	�,�p����#�>�aR�V����4�����ON���O�����&S��t)`����+e:�����p��矰�*T`�o���`N�pd������D�O
��>��Ɂ,Wr��y���?Y��J��R9e�Y��D��R�ɥr6�ȻB�'��%���'b�$�`��+%ʥ�.��UѺ�q�'�B�'����DX�tʩO���<#��@* h�w��)�.A-^���O4�Е's��''�A[/����HVS��d¡�����T��i���w�X�V�OLq�6�N�[�bDX�O�8	��Ȫ��{��O��$�Or�d�O�d=��s�ƅ ��X������?�2e��ȟ������D�<Y���� }� ��b�9@�A�ܽL�BH>����?ͧn `��4��$@�" 9q7��F^���A�#V�ęj����?�`�%���<ͧ�?	��?�ĠD��$,Q ň>4����"�B��?�����r}��')B�'[�S {��i�+� Lbd��D������O��D:��?� ���a���Сr	��h�G�g� ��/��i>�	�'T�Y'�dI��q5���1д�b
؟��	џx�	�b>�'�7O3s�m�󋒈%����?#9�<�����'��	ΟL%`�4Lh�K)Y�!�Шr2��ğh�	1��n�Y~�M��T�y�		�Z}�q�ABD�߬��5��	��<����?i��?9���?Q*�fA��C�Q�1��+@�-`�	p�(f}��'��'��O���yG��02��0��$Q��������<�X6M��|$�b>i3q���͓S`���uH؎P��s�B*`J8�Z���ص��O6�JN>�-O��D�O��S�� 'mx���[�nܪ���O���O��D�<	@W���	ğ��	
n�\d��	�9?S���R�-R�\��?y-O��l��?�J<YRLݳH�L�#fA6f�l�+���f~�G̠l!.�]���4���C�ӟ����'�2�Ƭ�0�p����Oд�{��'���'\��'��>��		A⎌�Q�I	I��k�aДjT�����D�O����OB��]�o�F�
7&(h��+�p����������u�hE禵�'�����B��?U��=�Dz7���i���'4�I�8�	���	� ��*�z�`0�S�X�E����g�F!�'���?a��?�I~��Lx$��8Bƾ<!�C$uo��(O�o��?iK<�|*�	��H�J�k�B�;9:��Cb�!A�.M PK�����-�0m���R昒O6˓�<�s�Қc��[vD��}�А{��?y���?���|�)O�=�''�3|c�lB��!*ޅ���c�2�'��O���?���Ms� �+az��#� 
bR^��fFU�[��ڴ������ ���l똓���� ������ 	�̐�S�?>���O����O����O:��"���ɼ���	
�%Z7$�e�L9�Iٟ��ɰ��4���d�O��Op����6
��%��[5l	j�ɩ�M�b�B  ��M��Ox��$�w�\��`kγH�mB�#P4�ح	�����O�˓�?����?Q�bX6��)O#'JJ�Ў-Ť����?Y(O04�'?��'�U>�g�_�-ނ9KQGJ?h�RL2��s�(��p~r�'㛆,+�T>��W��%,�Q&CB'8�4 �{O|�Pb�7e78\���T�ȟ����|Rnƒxu0�:'퇮ޘahw���@��'���'C���_���۴`R0��iL$qxu���׹:. ͓�?*O�O�<	2�i���I8*��]C��L1f�����pӸ)mZ]�T�m�p~�M�*��A�0f�剃E*ubփH�b#Y6]�C� �	gy�'���'�R�'dR[>)��C��:�f�P�`*G�=�3�"����OV�d�O���D�Ӽ��
$F ���l
T�� #� ��?a���S�'3`�\�޴�y�D��{ Fȅ�eJŎˁ�y�Ȁ�p�L�������O��d�:��K��/T����+ը^�L�D�O:���O���������������y�(�1��*�n��c�Q�	�<�''�7��ͦ�I<��i�>m�ܛu�X6T�nՊv`�q~r��l�ˤ䀇d�O���Ɇd��R�[o���v�Okp�؀��� _��'cR�'j��Ο�Rb霐-��iHUF�x00d"�����ON��<H>��Ӽ��KL	)��# �}V<�ʔ��<����?���P�`�hش��$�/�!��Ok��a��<�h=�s��;I�Mz �|bZ���	ߟ��I�@�	ПHi$f�Q)�PI�o��q(�)SEybD�>���?����䧏?)b���J0����E����5������O��D7��I�i�F���������E������{c�w�@=�'����n�Z?1H>y/O�4��d�(,˔فTēn��O����Ot���O�ɡ<��W���I���0�v��xR|����%>H(�'oɧ�\���ٴ{%�6�g�v`��]�N6θ���Ӊ	ߔ�;ӮJl*�6'?q¯_����	����'��;R��!�1 �Ofy��_�<���?���?!���?)��4J�*��#��r!ُTҤ������	��4�����O��O���P�^n/�����v�d�ҁ�_K�	�M�d���􄂘�Ms�O���T� "K�7`W�_��h��R�|�~�(��'@v�&���'�b�'�2�'���`�b� N5̡P�m�-&8��t�'pW����O����O����|Z2,��O�@�"��O��@E��_b~�U��۴5��xʟ"����Ѵ "}Qv@&"U`@��k��ě@"Ɨb	���|�C��O�%�N>9�͖���a L�,��㢡^��?Y��?!��?�|"*OJIn��~D��Z�CĈt����(�7Q��	럀�	����?�/O��o� b ��f���D�(�^$J�����tn�K6ZnZl~ ������_'��2w d�� h2q��	"|���	jy��'���'���'D�\>���JS��	�Ոϔ3^�x��E������O����Oʒ�����O�N	�p��"��0S?؀"�˾W��m��?	N<�|څ�X�Mc�'�d����R�����,�P �'��0(�	����|�Y������P��	di��Re�kn��h� Jğ�����d�I]y�>�*O4��ۡt�U�LP2m���a@���hO��8�'J.6M��%�� �$����".�@I�E��6A 5���)B����X�@���ڟ�r��/0�@b#T���!��k����I�@�I��G�d�'��iS֪߫r垽�b��{=ZmK��'�j��?���?y��w��
�$W�1��A���F1p���(�'��'7�րO ~�����,���!r4�$+T�oକ�� 69�6q`W��Q�"A&�|�'���'�2�'C��'*NMH��O;sc�#tl�)T��-��V��X�O\��?)���HE�%��5�'�T/8N�()T�S-�� �Ms�'����OJ{c%ػp�Kp��-�6���I�#󂁫�Q�H�PNN�K���D�	ay2�X�C�x`õ ��+�����¾+��'@��'��O�割����O�� ��]�7��������5�"A�43O��D(�Iyy�gfӢE�Iɦ��l%����aب���j�],@�lb~��Qk6,��(C �Od��1%�����U����%
�y�'�'"�'�r���:B^��q��W����������'���'�듖���O0�O��jG#��nE�[��%�ҩ+��&�<Pݴz��'`0\�޴����k4(q#7X2`R�a�2Wx�`g�S�I�v�Z����*b������@z��:��ԫ+�Y
b��y$@p��$Y�]����
�4]
����߳k2$��gV�[�h�r�&��pR�e�ߐH:H5��.ir�	�g�ԥGj��)� S�O���b�Ň�W�5��d
.)`���nH�7_v�B`ܱZC�����-ꮄ�3�,Z�M�F��8DT�amM�#wr����US' �#�Π$2Ы
%^��吶�] $ ��:5�� B�X	gO�Ub��Ŷ7E�q�R�/J�R �tn�u��a	Wc��\T$#���T�xX�ʒ�KM�����-�?�@�i�2�'[B�'�.��N�3&�L� %E�}$�ѳ;�d�O��|��㟠�'9�^���Ο��	�"+��h�oZ��$���T�ߴ�?����?���n��	�F�AC��1��V�L�?_&qߴ�?i��y���i��䓃�i�\��lU�Lcr�� �-Bj�	�M�����'��'a�,�>	,O�e�f�ܚ
��qnT71x��凚񦱢�E2��򉋯H���O��!E���g�̺�*�&�Aa�����Iٟ���ğ̢�O���?��'���I� �9dt���g���l�"Pێ}�6�y��޼�y��' �'fh(S�ʐP�6��CF�[��%��nwӨ���OX��'��I�<&�֘�T��G
�uČy1��/N���m�^���?a���?J?A�J��*l�U�V�Z�g���W�`�Ф�'�	�,%���I�@���w�@�aH�PG�a����.OV����;�x�	ʟ�I֟�$?M�O����֯��"�0R��ͻBw,X�ߴ���O���?9��?�W/���$�����Ȝ�;h�8Q��YM~�ܟ���ٟ�`J|�EW?��I�}^y㠅	6Xv-X���cG��ٴ�?�O>I��?1��G$��'����e,W�7�Q�C
��SN̦M�I꟨��g�H�	"����O�D�O���Î�O���	��ҝt��0{P�MP��埰�I8[dhi�?i�O~];]	tB��Ŏʫ]�`�شx>]��?a��i9��'8��'�v�xZ,�c.M��½�&��&]�>��G�itb�'?����d�|�O��U9�'T�Y\Z��˄$tS�=j�
bӜ���˦��՟����h�O�ʓ'��cP/B�?� ��M�`/�8�a�i?����|����<q�/�2D���'�%Ƙ��9i�I��M���?y��?��\�L�'Ob�Oܥa$��C� ���e4RL���ğ6m"�dN�X���O��d�O��s.$cx�Q
���30[�<�1�榁��ݟ\c�O�ʓ�?�O>��)��t��m��E�v|���?PBr��'[<욄�'�|�'C��'�~*��B�լ���'݃���7��٦u�O�˓�?�O>I��?)#��+%����ϓ�T�Ź��2F�{�5̓�?9���?�L~�0���ô��"��!a5��A�H��X�P�	�� &�T�����'����U�ݥ4��cՃ�n?�1�jU�y"�'jR�'^�����O_r��^�����åh���;�ȟ�^�6��O֒O���|j����3��UW�ǶD ���;6J`7��O����*N�d�O�t�O��'Zc<<� &\��L�)���4_d�YH<+O��d�O|�����P��F̊p�����㑜M�(���i�$u��'��cp�~���M��?���\hd�:N��Ń4�RW��T2�o}����?a��h�O@�S
��6I �t�JRKS[���LK�k}�	ǟ ������џt���� �t� �ڵa�#Z�4M��	�,.\�'��,���4�ʰZ�������Bf�"���K9��A%`ߙ�M3���?��?1+O��^�� �5M|}�s�G�[}V�Hb��8c�MDx�s�Q�<?����?�;-0�1XOδCǀ�qU�WF�Hn�����IpyBD�~���<®�y�Í72�:)�HX�|�O����	N�	ܟ��i>�x�8]#v yt�r� 0���mZgyb�'0��$�O����4m �N_�Ao`�*c	�C�6�Lr�$p×����֟�[ybПr��"i��Y+��r�jL�ub����i@��'��Ot�ĵ<yB�Ц!RbdǔA���ƃN�K!x��Eʝ�y2�'jB�'�Z����O�rdG4h��;�A�
tr���e�ԋ2;�7��O<�Ot��|������E"����� 7�Z}�)O$6�7��O��$�p6˓��i�O0��Ok� ~M
�g	,i�$�0r�	6s�X�b�xr�'��'B��"<�;_�T��c �kQ�x�s�37�)o�#����ٟ�y޴�?����?9��J����m��̪��Q2]�ba��ؐ`|V7��<���?����T[>�R�d�jѐ��r��c)E>5�a��i��B~�`�d�O���O��'��'EZt�ѓ@%+��r�O��g��DmZΟ0��֟,&���=��b�����5(3�IyCHA�)�R|�úi8��'y2�'|�)�J�x��(	j����N�m?��Q��N��O�$��9n����?1���?i�wa J��w|M��#V"x`z�	��i���'v~O�S]�	>P�F�k?q�N����,?��*J<Y�i�����?���?aI?%"&N�Hވ	�GߵE�X���*{�D&���I��$$�Ԗ�uGL�Dt�)3� 	�<��c�J%�MC��[��%��?����?IJ~�S=�$x�ufU45>nIX�۽lv9�ƺi��⟈�'���'�b`�?���^w��q6�S$%�@��@��Laz���?���?1����'Q���۟�X+����%�ګ9�%�g6J�^6��OB˓�?���?�����<����~ҀD(	$P�sIωg|�RP-�M��?�c��<i��PS�S����I��d��iA�wƂ�5�[��<���$�OX���O�iS4O�ʓ�?	�O{�`Cn�z%DT�2JV����4S�6���?q��i���'���'VX�Ӻ�R�EA޸�n�=n��p�$E�禽��۟��gc|�l����|jƕ޺� �bk�����G=s%P�9�N��E�ɯ�M;��?���?9bS���'�p����j�T���z~����fs��9�7���'��' ��՟�z���+9t��P㐩T7V0rh�2�M;��?9��?�Y���'��O$a�u%��#�2���jN8��"��7!K�d*G-��O����Oz]�$6P��Uꢌ<XTx{�L榡�	Ꟑ��O˓�?�)O��ƞl5�� �ء2&#*y"��Y�i�⬏!�yR���L���'��'����5�AH#FA���f�	/֡��
�M��X�@�'IbV�D�Iڟ ���<u&ӱV���C�d���(e���n���Bg����	ϟ����?�O�6�6P ��T�������..6�<�����$�O����O�ȇ4O����<sz k��=S9~�2!E)G����O"��O�i�;��L}����5��;���0��n]�QI���M{�����O���O�ɛr3O��d�����N�#���q������)s�����O�	��<OJ��@~�t�'�R�'��EX��D�М�#����3ɴ>���?Y�e��Γ�?�)O �(y�iJ#G�^	���i��6�07�P�2���O�`l���<��ܟ@�ɥ�����!��]x�`��A�D �t("�i��'�~�[�'@��<�.�t�IĻ�tpT�`���ұĽ��ۥ�M�����'�b�'y���>y-O0�y6��NY�ID&KM�y��h�٦=c`+?�.O��'K���Χ�?q�E r��њ0F�HTd�q� [�`g���'�'N���>�(O^�D��+���S����MV#@2���"�>�,O�h��9O�Dx�5���$�O�D�;H-����±Kt�l�h�X�oZ՟��	?���<�������Ok�G#�ɣ0 �4lq>E�ׇI�Uz��
.���IA�L���ߟ��I����s���	���r��uT���cB�^��6-{}�U����xy��''��'���&!��E�D��JI�	���yb��+1U2�'s2�'��TU>%;�O:��Ja�T<,f2��FA�,Y6ms�4���O@˓�?����?���w}�`ÙE�� ���aT����ʚ0�������	ן0�L|B \?���E?&-��*�������4L��4�?�.O��d�OV�6w�i>7-�S�hS��Z4!"��b�MJD�f�'8«[,�y��'N��'�?i���?��.�0K�Li�#�"��A�A6<�	����ȟ���O3��4�"!��<���c�i�PJܩ�M�ӫ�<!��f�F�'}��'DR��>��yX��aRE�\��g�h̒�m�ן���#[����|�e���+��އ-"5�P���B�f�{��V¦=�I�M����?����?)�T�̖'�>�jч]
&<@���.,n�	���`�R�7O���<�+�.*r:����� P�	��Q��i���N#R� ylZ������P�	�����<����~�+�� 0tL�m��\��ՒT�����D�<�B��<I��Y�|b��?Y��[81�T�
U&l
QhJ�{B\ҵi���'�들�d�O���?�1.8�L+�B@\X=���a���'�p܃�'8�� ��'xB�'�b��yZw�<(�r,��V5@�{s��m,��4y_�I}yb�'��	�������l` ɒ"[?$ŀB�B�(; ��s����,.���������4%?� �O��X0��n���b]͔a�޴��d�O���?���?�0���<!���#3OƠ�`F�TgX��s+�y�����?����?i`����~*��3Oz��f��,w�HT��+)Sb�궳i��T�L�	���I�վ�IT�ܴc�-93&B�$3���a"P<hz�lZ����.²�	���A��f��O����a/Hy���6a� �$F�R�]�'�"�'0��/�y]>�b�7��mO�U��k�<H T����릡Cv�(�	=�M���?	��?aP]�֝5�����ע*��M�C�
U07-�O���VD�Df��'��Ӻ3�*ם_�ڡ�U5!������~��6��Or�n�������I���<q�� H쑣��I�
h�1O.2S~-���i�a�'<RV�ĕO��;�O�F��QmjP�)T���0�M]7��O0���Oz�a}Y�p��|?��H�9E�Q�c�2��Q��@Uڦ)�	��l�� am��I?uh�ڟd�	��8�FC;���{r�Z6u*r5�Ɲ�Mc���?	�^���'�"S���i�mH�̚�=^��R�?�8*��>��e��<�3����?I��?y����Ӻ��f43Q�a�B�7J"���U��m��}��'J�'��'�^�@E*�Gx��G��(�`�*\�ў'���+�'���'�R��$(y>�Г��
���@��L�.[�=��>9���?QJ>1��?q�I��?�G��-�H��.�( ��({���
⮔͓�?����?�֑��ΰ~���/�f=`s��>Q���ץ�!�ԫs�i2�|B�'�N�#�y"�>��ˁ(�����Y-	��a�X��7��O����vT�d�On�O1b�'C����G ��_-n]|x�㢒��(O����O��;�+�O�O���1f$d� �J�?i$����^�6m_;S���OV0n�ן���ş0�ɴ��dٴU�H�A�_-M��t.�}|���'�⣖�H���|�Y>D�eӔ��"kҜ�R� ���p��i_B�aӪ�d�O����O�8�>�"kG�m���B��P� �@y��G>;��G�x�R�|�]>�c��u���I$|���W�J��ջuE�<=ݨ���4�?����?��8�'�2�'��*X{�ȱW'��~�"�Y�@�g̱O@��:O���8O��$�O��$�KhT���oV(�a�ʁS`�n�˟P�ɴ�ē�?�����2�>?���qjfr���u�g}R��U�r(��y��'�B�'y�'\�Ra&\%X3���1h�0et�QnZ��'��|��'��H(H����c
��|���"I�H�J,Cw�'^NA�',��'�����d>�Hug�#��h�gC#%�8��>1���?�I>9��?�Adڝ�?�3��quJU�G�B����@����q�����?Y��?頕��N�~��quTtcD�	�>ђ���h3���1�i�|��'�"%[0A�2�>qŭB2E ܨ�0#E�x5����)�Ϧa�Iԟ\��@y�X�I?����O����O
$k���@PAmJ*,����dDJ}�'R��'-T��S>������`%z`��*�-�XP t̕��Ms�C��<���[��&�'���'�0?)��Yj{��$!�I���(�Ȧ9�	ٟ��q�%� �O���!ܴYeX$+�/�����99�MlZƟ$�ش�?!���?���p����!LRxp�PΊ-Tԩ��iY ��?I��O��)R�'l����6*�p��odx�C�\�7��O����O����s�i>��O�uY� ڭ4���!o��[��5X��i��O���ƼH�D�O�D�O�18��L++O�ٛ�;Os�4������쟨�'zh��?�O>9�Jϝ+䵩�CԂ4�ŢS6j��'�Е1�e��y��'���'��s�����=�ّ�%G�g��m���ē�?I���?!*Otʓi�����N�)n��D��_�T��E�<a���<���?����,�j�S-�(!�/ƴ�p��itOB7m�<������?�,O`yQ��i�� G�]	�e$�X+v�<b&�������I��ħ8��ޟ� �,��j��4���
���9�MK����?A��1^���>i(W45��%BK��Iq$�尿�	៤H��v���	���	�O��$�O`y�ʛ�a�B��L�fπlQ�.k������)��#<��OS0���
G��Zl{�o��)�h�ܴ ��ϓ�?A�iz�'���'�� h4%AŦ`L�Il9H!ߴ�?Y�Q���Exʟnt�w�i̶����Z�n�9F�h�hD%NЦ��	��M����?���?�@�d�ebpD��xO��D�Srp�l�w[0"<A,��{;O��ė�&��li@��%3���Hl�������I���'&"�OX�M�T�mI�
5D`�}���$�?A�ߑK��$�OB�D�O���O�]m&�i3��GU���A�Qݦ������J�}"�'�ɧ5�	�$V��`����x�Xh �P���V/�~�Oޗ�y��'�b�'�'4�zZ���0��ܑD�ρW�oZ���'�b�|��'��-kɲU�v� (bn|�3��)Pɓ�'H��{�'��'�b���ou>	Z��V~*lpX ��	x�I����>A���?AK>I��?Q���e}hȐ1�؀uBY� ���'^~x��ݟx�Iȟ�ZwB��՟��ٟӈ�1���b��%����M�M;�����?1-O�,;בxR)�8
��Je���t]�4'b��M����?�bAT�<q��]s�Sן8����G	W|�1��E�|�D=2&n� �M+)O�ʓ5Bl���🛶�'tŸp��v~6L 6,�$�MsA��?I��?���?	���?A��?s��3~��hSa�{�H4��I/H0�f�'l�ɨ��"<ͧ7�v�o�L�D�c��I<BHE��j�F.V6M�O0���OL���OT�D�<�O�D}X���&.e��#㞒]fyzb�>Ѥ@[a����A-�y��'j����\�=�~��䜆k�*	���m���D�O����O
�%�$����T����E��>O��D#d�	#"A �E~�X��yB�'o2�'�~܂�o�%@�X�P*�.\���9E,o�����O�H&����ß8%��8� �uر�$X8��b
�3MN ��W����g�d���v���֟\��Y��@#.,@��ͅ@N�r�̽T��F�"�d�O���6�D�O��d����S�@2`+��3� �d�I ;O:��A=O����O0�d���ʧ�?��ϓ-"V|	��8,� ��tnБae���'���'��'��S���&Ӱa���ϧ
T�%a&�	?��������<Q���?��`�O$b꧅?����d*n�9�)
3�Y�l�=I���'4rV�ܔ'C���ɟ�	�����uɃ�[��mQ�%Ӂ5�Z6m�O����RU��d�O����O����O6�$1be�uA��
�쳤#�HA,-'��	ny�@��O�nZ6\Z��U�ܖ'������u˛fD���y��'�d6��O��d�O���NL~�Mؗ\�`U�v�_�p%�p�@L̮�M���?Ԭ�J�'��#z6m��S�����j�T��`śv�'��7�O����O��p�s�<=��"�hը�I�D�M��iż���D�|j���<��`.���s��!{��CP.*ohZ�i4"�'"�'�&O�d�O���:#C4�ٕ�(���H
V��b�$Slu��*ǉh���I埈��DV��)o�`l �A5L��M���?�5���OV�Ok�'4�5PB�P�j��H��D?&��� $&��	/��IԟP�	�X��.�� �+}bfP�'����Q�A�i�&���D�O�˓�?����?a��3�D���T�::���d)�V5ΓL��Γ�?����?9K~"F0���qE�1T*(�P�M�&{����i5�Iݟx�'4"�'t2a�.�y2�ʡzK2 `DjC(.��@�>p`�Q�'�B�'C��)��XC�D�'J2�	0S=Y�n򧞱nޖ(i��f�D�$�<����?��
����ܴP���Qh�#�,�%���ǿi�'�~C�'�Ҫ�~j���?���*��PH�/$eS�-�H�ZA�T�|��ڟD�I�]n��d�?9����%�}@��-l[ ܡ�f�F;O@������IڟP�	�@ �O���f1fűb�Q �~="3.�==���'W��]��yҗ|P>�"fӬ\X�HL{�\�`�\*�@Zr�i��oӠ��O��D�O���'���4p}���6FĶ, J�(��$ƈ�:ش<?�a�����雾�����g��)�ӫ���y�e���n��2�� �KbH`)1B�>Oܾ��R�������7�Sk���Rг�銫Q�ɠs���Y�Ƚó�
:e�����,pH:��4"O�p�wꍥM��)`򀄣Mژ[abA�L�(����yb��X���w8IR���;� i:f�M��$�y1�)#6������mJ�Dq� �!/�)�!���ХP�
S�d�Fy�%�L�	13~z�	D+^?v�T8rq�
w؁�F"��J�ʅ��Ȇ&S�УƯZw�gm��
��Y-&>dHC�۰,G����O|��<����?�OI�����N�jpC�l�+i��� ��Y�W@Ȓw,���k�� ���a����Tg�'�|ظd��* 4�#DM��}a{"e���?a�?(|̛�b�:F�� � ��e�8]P���)�|d2]#��&"������L V��ȓ����&��E�D	�J�A�����	cy��Ѽo"���?�,�Ьk3���V���ᖄ�$J�}[A<O����OX���#"�0j�F�`�O�]�f�`�N2*%���@>I)^�<fd[�j�&9*c*Dq�<	��L�
��4�@L�FVf02D�ɢB4H���O��?��aƦMe��K�J,lm��a�t��I��,)#�%WO��0�;M8��d≕X��1X'��3�0�萫F���?m�;�O��#���ON���O�P[����8Ǹ	�Uξ����/!����pN�J}*hJ�F��ʧ��?�b��7J�A�
}a ,F�&w�H�bMӪ~���p�Y+���񧈟2�05i���sl҂p I{��Js2S��'�"�����O"��#�y�Y�$��",�x�sA"O6|c���6��@�a��${��"���HO�өj����A�)%ƨ�Dˣ������)�o��M����?������O~�d��*������P)2lx�HbGL-P���ߎ�)`2�K����I�%��5P%[�H����N��E ���^������f��;ǓP���s �7��A��ڼi��T� sH �����G{^�$��N՘vN|�z����X�".D���B؃td� �N.P4쬡!J��HO�M��3��=�v���E͂��&��ͅ��d���Z���NX $��R�$���jYw$\
t�N�2h�̆�@Yb4[ɓ6�1����k^h�ȓ*2���w$F�a��I&@�����d�-ӕ�=xF�y(;H��ȓ(s��c���R%Jc�� ����Z��E�P�MX�"5�9#]�0��MWB�2Q�3��e�v�C�1�Ll�ȓ$#�u)E�+%i.\q0)�PZ�!��S�? �}�ǂ�z�@��B�	G�<��"OH����H���J$��3\��"O0�+�ăL�\�QT`�:@S��"O���U%=9�0D�6�DWU0U��"Oȡ�/O�XQ6��3E�$�H��"O0!Rc
��^�sD�8$y���"O�kw���m�L �C��k���2"O4���m�+#�l����{\0Q�"O�`�f0)a
�"r'�.kTy��"O�T�R-_4B&M2Q$�Ksʡ�#"O0� �I\�q�y��M	Ok��I�"O�|�E!�n?z���(�#j`��"Ot��	N��XQY-x�"O,����=k|@q�G&�	����"OA�$��6D؀��0��T��bQ"O�ؚ���bߜ=+�b^�8J��v"O�Q�fl�4�HY�uk�s;���P"O�u�Ba�G�� �$�1-F[�"O�5��	�&UR��D�̍ˡ"O���ˊ3	'T�	'"D:V�-�"O~��H�N���C�ܫ< p�1"Ozr��/Xx�}�w쒒&(��y�"O���ǥf��{��"��0�"OHi���̗�.d���k�F|C�"O�e�&G	 =|�;����k��5�&"OT��V�Z�yH��2Ԧ�r����"Ovx1bN�wHfI�#d�o�||ؔ"O���c_�X��ɒ"I��
<�C"O`ii�f�F���e��"��,�2"O���B�6�����I0h��yP�"O�}���r�����݈c���#�"Oj����=e�(�0gҭ=�$��7"O:���o� �S�X��PU"O����۲AcT�q��g��!"O���E���o(eᔣ�mnp���"O�I1D�;a����́1<��Q�"O,�[�fό/��'+m��yA�"Op���i<x��Ui�j������
O�Y��CV�n�>�ce)�W�t%�W�2t��#�^$�M�%)�.���k�`����	6����{�H[�N9�8!�!S�W�ye��4�yRAZ�.���F�8Î�ꃆ����It0�=ɍ}��@J�z���(�j� L�.�y�@)��(ꔡ��T����Ыی��'O�T�Um'O Y�G۫9	���Ǌ] (M�
O����<=B5�j��N	A��7>�\���}Ȕ���W98�H,�*�[qN��	Z��(b�{�ύ,:</���1��ȞX��EX�'GV���� �lUQp#L�8�Ν�N���"�G��ا�O���2�nU7#���lߍ-�	)�'8J�a5�A�k�.����L�}��{҄�"����dP<F�H�d��Gm��0��&O̡�$�g�ТL��4����\� ��U� o(<�剤����F�=|�l҅�Lj8���#���'�>�'a�-q�V�'�H�5A�5��'�v��6HO�_�Xs�Β(1<�XL���f���اu�{�
hM�p
�-Ҫ�R�L���yn�:Y�*uH�EH>��X�+T-��'�x">+U/�y"���Āh$��<�^��)N9��xB� �h���@�d_�6XJ�5S# �\�=1+[=��O�!�%�ߙ=����P��!&1�hc"Ovu�/��(x-(4(�b�h��'���� �'���G�D�xƘ�7�Y%=T|P�u[�u�O�� �-1��i8�m�O"(1�"O� X�F�f3L�YfL�z����C0����$�T�d�W�9�`�k&b��n]!��3-��,�g*��$�tH�!�7-����)��<S��K����S��J4��F�`�<���ʉd�����O��;�(�_�<�ꓛh(p "5� �Rl��MR�<AE��9-��(%k�$N6�rqO�<�!�*�Ԍ0p̉�u&�&�Ay���3#�a|�"\�Ws��[R�En͞��D���>�vD��yb �a�q���ZY�8󒦙�y�%�Mo�U�T�b�R�����hO�Q�&D2�'�@ ��[j�d�1K�S�XĆ�[�U���m��9��
-^�I,2 ��?E�T�A�h�����o���l��I,!��/A�(mIp��HZ�\��K��;�ɇ20I��I�����ČK�2X��ѓd�>B�=F�>�Yr�֛��rJ�K B䉐"��!w/������%�mp�C�o��%��J�"�^t�R�M�P��C�	�wi
�J
�|*|`��̯
��C�I�[��8ԤXT\$Q"(�u�C�2u��t��׬s}R��D��%D�B�I("�F�x�
,8Z�I��F5k$�B�I��
�8E$��*L�ir��'g��B�I��Q��/�/3xDa"�e�y��C�	m���w(A�A��("�X�!M�C�l7]!P R(\z�x��C�	6E�@Sq�Q�v�p�ӫe�*C�	tcMt�:nކ0��	S��B�I4��w�ʝe1��4��`��B�Ɍ|�4��Hx��	�!	Χd�B�I	Ht9C�χ�nP*A{�j��BB��/L�6U�#��<�V|�t�HhTC�	oPx	zE ��):�m�e#��8C�I,�F�r�m@�������X5C�I�3]|Ax�	P$$Ш�Z@�պC�ɱx�t]S�*��
C�yC����.+�B�	o;v���ٰ.s,`v�Ѩ7��B䉀/`���,V�h���`�(��^�|��������3Ѫ�(�M�ȓ91�mˣ另G��Q�S�/ 8]�����X�
�> �ܨBJ�6|f�4�ȓh�����o��r��s(�4o���ȓV�(u��׻f���j%߸Cј1E}�S%=Yj�+��]���Xs�QY�D�	5�F�"BNX/2HQ%��b�NY-6Xc��>�8R��E2lrT"� 
���E���`�����@��<?E��K��*�J�m�Pf��7j΢�Y�I>Y�jϠ�����!o
Rf���o25r���O��]�'�:D*d�.A�U���O� R��!]�4���őjIJ��$�x8�H2\O��Þwt����_�"��B�K�Ƅ���N<8<�u��f�7M�#e<���O̩�&��W�~Ũ�AA D�ؘ�5�ɞnc��;��V�^��F���K9
K`�SЫ
�3"٘�����'�G&o�d�!0��FW�S�~2hT��F�3�J���8���I'<B�	��E$"h��S�84v4���G-_e�,����u��0	[�6������؀(�� e�m�ܳ��O�Ÿ�@�-���i�$�� ��	�jMr� $Ć��5{z����' &*��#c�5PL�(r�Bc��q�Ә?:vxC���Y1 ��>��M��X/R=\<nZ��QğI��A�O�IVT�6h"Ο�hQ_:����G�����o��y�L�?"9�N�?�D��7G�c�̕�'��`P��7D�:�`��["M���)��f m "�ҲmيqC��D�	��z�dK�"\!(Ui��xZJ��r
M L\�q�c0kҠl+�̀j�qO����fAw�g�$�g�m��_�_�4M
p�B�&�qO&�R)V3?ٴ9�f˘�c?���5vU��)�F�y��
�˝<n��}#��hc �+Y?ML$�$' *,�x��2�!A;�����T�	��l��H��)� "M��lZ������k�=49�q"f"O<�"�K��Zx����A�9��`� �i�z��R�r�>�8�4L����M�ch��X��\�u�J�g��?y��{��;֜��C�]�#���A����}�Z蔎�,%�p���<�Px�h�_|����G,>;��������9E@L�烟#z���?���k޵[�h �F,)� �˱�7D�d c�Ր�,<��a��̭�'��OZk���3>��i&�"~�[���	!���0e��y��KD"O>�p�+Q��Y�QҨ�U"Or,��� � ���Z�6Ȥ��""O�x3%ƛ*$Q~�kf�ũN�� �d"O�|�M�6[p�	�*�k�l9�`"O�i Վվ2,�m	�e���ö"O\!S��(tX�A�An�l�G"O�y0�͐�v�\|wT>\�!"Ofx(�b��;��9�oZ$*щ�"O���,X#I� �r6NѣF�P�U"O�X�a{������O�& ;r"O����׭.
4B�iF�L�d<9�"OF�b�nz�Rɸ��Pw�|Ȃ"OVa�FI�o����׎��@���f"O ��T��$'V��:r�/d1,�"OZY�Ѥ@�_Z¬×�!&��i�"O���� -p\Z��TQ,Q�R ��"O�0�e�G�&�4��A�!]t���`"O���R��ʲ�H�!˷H?�\��"O����>AHdȔ���&�=1�"O3���M˲�(�Fԫ�h)��"Ot�����ۮpSD ��Zþ@x2"O�Y���J�t��!p�DS�AS��hF"O*���!$���aUCJ�f�Ni�"O�da���@�L�03��4�f@�s"OVA��
E������Jl�Ԩ "O��t�� I��W��	?�v��a"O�d�d&�s�T  3�~��"O�p��ױ�� ɦ�_�g$��+s"O�`�VΌ�1�^5�BD�5f@��"OL�`wM��^�HK��Yi��q�"O�a�!�&����+�R��3�"O\�ڒ��8)-�"�'���c�"OXYA��[���LOD1x���k�"O�u�q�� �E��M!g�\X"O4]HfiA�^궵!5��"3v ��"O�5A�ΩK$�p���\�x��"O���+�lS����t��"Ob����&*�ެz*�.W1ʳ"O�T 5�q 5�H�s�Za�w"O�`�u�
%yἼx�GO�YB���"O��{�JR :�ȝHtF�+�\� "Oh�a�C��U(pFY�<z��"O��x��	�>�P*1�Fm<<��"O��S�Jd6%�U�OqN6m��"Oz��b�
L��p͎
3B��6"O���F�,�|���̅��؛�"O������Pt���we�8p�� �"O|��H�{���6���g��z�"OjIN.S�l���` D��6"O0(�D�P��]����@��I�"Or4�4��'2i��O���"O�P��ޅ/��%z0`��N���"O��
��L�Τz���)^0(�"O� ���{���˷hǳ	ԂT��"OBY+��7��5��F¡63Pܠ�"Ot,�c�!jTJ,㥝���q��"O� �|B4�ǄE�ؘ2eJ�G���"O:��v
R�
tmC�4$�B�`�"O<4Q&F�U��Q�gN.Iz1"O�MaW��c:����+��Q��"O`�IPJ#|e$@�0��LS!"O UK���2n��[rK�� ���Z�"O���#���:�6�*�7 �#0"O^���L΃} cq#��B�� �"O��!eI��;g@��#K���[�"O���A�ܠ\����ADh��P�"O�8k �J�|���rւZ����ia"O�Թ&	�.�V��T�B�+U"O֡p����AR� �#$$��"OhD)�"�3����b@��Y�̼!�"O�p��e��.>�0h��';쮹�"O�ԁq��u���m�q�^A $�'D����Jٰd�����6ihn&D�$;���&e�)�G��*3�Ν[��/D�|�V�Z�zQ��Ӧ
~�iY':D��!2�Z2d��W&E�A=`��<D�8[ ׀F<�d�W�a>�AB6D�dґ�I����7�AR* 	�S�9D�h�F�W�~0�F�I6��SW#D��)�D��(�h�m�Pj���#D��4Hլ<�l��A��|22B4T�$ �
��(KoC����"OrU��ݦt%����"\��\x�"Op��1J��'z���Ơ_�R��"OV좤�	���AR�v�YC"O�U���)�����?C�hL[�"Orx d�"�q�]�L�葙�"O(x���F?jl����
=%̚u��"Ot(X
�	1��H� D�`"�yK'"O�IӃ[3<��M�`�P%^A�z'"OT�*Ā�:[�����>���"O~�SCL4R�� �����!��&"O��"��7^��d`���e�dܺ"OְZ�FЦ���@�Z��b"O�ᐅX�`�с6��_����p"O*�R/ʳ#}\$J���&�05"OlT��b:p���!��A�/����"O>�s��ƃE��9btA&3o�U@�"O��R')�Ƽ��Ù2K~�bS"O��;���c*f����D/c6�+u"OZ�d���]�`�9dInP
R"O�4�DµX��p%X>u3�P��"OF,��`�@�P1&���<*l���"Oqs f�F�l@�c逵&9�#"O¼s`*F)ch ���- �"%"O*p��J��I�f�2^��a�����		{�4�UJ_����J��{I\B�	�n&8� T4�8b�^#;�C��):�4����! q�����DFvB�I����Ũ�?�v����ƶA��B��k0��B&�A%+�t��a��3�B�ɦZŰ� fJT.SDu��,se�B�I6bc����G��aB5�ċi*B�	+kf5BR O��˓f�44�*B䉣Q=tmXe��|�aZg���C�I�f��Tȑ���gyrA�v�	�v��B�	�Dh�<�7m��i7Jq��IS�rT�B�I2�~�yԙY)��eO46ϞB�	-I�6����@
&B���{QtB�	�j6�6'F(6����oS!`�NB�)� �%z�I�{�M[��]���B�"OxI����LӀ �7�7�*K�"O� RcU�zeZ(qf�1��R�"Oz��d��-P5@�$J�>9��"O:�ãO٤M����V�Q4o�t�i�"ObPrfcx��'$�y����"OB��vO��N=:��e/�a�"Oz�A')
h�Yb`A��)�@�"Ox%��mթ^(�rG�x�Y�"O�,��)J۸�Jd�^�2���r"Of��ŤWc�i91�Q-y��u"OJ8�0!	`e6�Y���!c���G"O��Za�I�	 R�J� ��e+�0I�"O,���f�
 �̅Q ؈w���:�"O,��N�����k̖�6,���yr!�(}�� ��U�5,l��&A��y�DL;=���j��KVU�4pw!�'6]���3BB�����,��܊�'xDP3����P����.�+���ʓق5���S2	�h��G�<c���ȓBn��銉5�:h"iR�3�^���m������(fp�1DM21��E��l�B<�MM;36q02�O,Vh����.[�*WR%~���PȨ=n���ȓ�H��� �|���qFg���XՇȓ��x2�i����ă6]n@�ȓ}��a��'I�Z�Y��ɳ�4Y��#�&8�&�4��퓒��J����=�	�.������J_$t�q��0z����ȓ��H�B@�~���y�/ƪ	�Іȓ��D b]��	��������ȓ�"�*U�_9"u��FI�5�d��ȓ �8s�+��[�}��'�|+Vن�Wx��1�N�nT ��@-���@���F�p�!�����N)H�<��ȓR�J�UoD0T(��R#)>n��'_`�p�"AtF�"V����Շȓ_�D��A�#:��d�`i�4����>�����T�xH�eMΛN����JO/�y���9Nr��sl�@z�T�f��yb��*-9%�,H���僬�y�a׿j_�أ�j�
Q���X����y�%Hrd-P� 
]}l�2���y���b�i�GHI�UҠ��G�J��yrE�8e$� �RQYҴ��y�K�;1Ԁ)Ս7��lq1�Ě�y�� \j��r	�v#��f���y"-��q�X���͔#,4� �
Y��y�ޗ[�VA�BE�(�j��A@��yW�b�FV.��#t\��	� �y�J��x��ä�8Lݪи�M���y���~�Bt��Q��h��G��y"�
�K�LU!If�	�)�9�yA�1T<��ɉHgv%�#M�"�y�揣6��t��<�;�bX�yY=({�	8���^�T���F��y� �qN\Ѓ��W�� �����yr���x)�m0��"F����DaC	�y���zN�u�ӋχC��j�gW��y�d�<z���q��X#;1�3�Ó�y�Jic �X3FW�^�	�+�.>��|��	6W��ug	��Mq�E�NQ�s��C�I�$��p��#ǜ����ԾXpC��p6Q��Ԁdj�uN�C�C�)� �ղW�D�L	~�p�(׋Fm��:�"O����"[�:��p�d�}S�q�4"O�ub��/#�A��oX�g��tR5"O�qaB��r�2�B2H��e���2R"Ou3�↥�ݺ�g@�z���"O��Pc��j����%.Y�B!��"OZ����Øn,I��"ƫ%��͑#"O P!cN��Ry2A���J�l��U"O�I��
8 	Ԁp�-��1H�"OA�� %��-T�/0h3�"O�L�4s����鉱@�`�#�Q�<�q�׼T�n�k)Ϫ���t"؄ȓ3�~I����$r�X#��>R셄�v�%r�ϔu)��އEm����&\��V�$y�(��Y��ԇ�ͥKz�ʔ ,��d��U�=D�@0V�J�TnN�B�]�]��=D� 5��1�e܆�K�j:D��ɣ��3(��a�A�b��x�'H�R��{"�y���;Z"^���'�(J�h.g�VL�N��:�� �'|�y�'�:JI d�D�[�$��'(���#e�w��La�*�gRN�	�'&8�Δ���-�[!Z���C{�<����!�����*��a�@P�<9�hE*;F���2�
l�XA&�UN�<1���$`�4�xC���%�nt'�K�<Q�"]<cv`�����J�V��% I�<���-��8��É$��dab m�<��Ɣ;'2���/D?p��e��f�<QC+�yH�#W옪�te�%
�a�<���(V6�#M
�uX�d���i�<Q��R��-�Z
�T�N�::�C�;s5�1��e�	
�a`Y�C䉃G��ypc�x_���b�����C�I� ��+v	)�X8k#T�|�zC�w���N�Nd9(q��e�<C�%�2L�dY�5��܀R$D=\�lC�I�'���N�q�X�)hB�\9�C�	�v��PD�kՆ�� l�:C�I�fq�ɳ�%�9C�Z��*��<�XB䉷>����E�@��@6l[f�C�#V,���)V�T��	��`M?3�B�3G �@�S$Ə-���s�4c6ZB䉔'j(��0J-[���a!?y8B��^��zff%�ܙKB���B�I�Y
��u�	 �~��M <~�B�I�'�}�ծ�e��`��k+U��B�	������I�| B����B�IB��DJ�J�-8�`%ҹ<'�B�	g�|��a	ǘ9�쩺tot�6B�Ʌ/Q(�Ȗ��82�ٸ׎�>2B�	#H�(!` I��T��rb��l"B䉌%��3��'%<��$@9DK�C�IN熩Y4b�d2@`ؖMtC�I!8�u� jd�K!��OI�C�9X�E!֡�'0x��nM;4(�C�	���\KU�&yGB��c�2N�C�Ɋ������eP�+�,��hz�C�	�RO䑑��i���!s
QKDC�I�D �!�����1(Ә>�(C�I
P\�ħH�a�o�4C�ɾ}�}f�˓H��ÑL'm#�B�	A�(��q�%u��Xd��y:�B�)� �ѱ䎊>s�F�R�N�I&R�9�"Oة��;?`ب۵�](���"Oxuo�LW�c��?7�u�"O�H`B �/TP��B�D��U��)"O�$��TJ�fI_%N�(!4"O,H���xٰ1� #�Q�"On��'i�2K�� �A�Ew�T26"OeEȃ�J�j�����b
���"O6��H��*� 1�!�0D��s"O�M��M^
 �eZaGY8Q�i&"Ot��f L�K��b@�Z�j�fX"�"O�m�W,��82np�F��K�Zi��"O 4 ঐ0ܲ1�&_��F���"O�b�z���ӥk̈���"Oz1h�&��K�.eqUkͮ$,h��"OE3��$):�$H��^�q�(d��"O�t����
O"9�tP9\��Tj2"O$��6��<w���J�MUsJ�["ON�j�园BPj�*6"�l3l���"ONX��/�.l���!�GG(&���"O�YSiΠZ����ƒaFn��"O�M��H�&?@(��˴�0I`�"O��w���P ���r��7"O�!j�i�~|ʼ!��ޣF}41�"O������$j�XAŔ�bF�y��"O��A���&���B�ʰ1�A�	�'���Fȷ;d����ℓ�L0�'�d�8SK�,lfH9�)Y�w�┠�'mz�AA)=QEM� �Ϯg��Q��'�L	`�C�U�\05�Z.����'nD@�vW;�����Y͆���'�ĄQ$�Y){�H����T/.���'
�0
r��MIT�ˡR$�yb�}h�p�&C%:W������/�yMW�.y��+82̠8!(K��y���SX�ဎ�'<�X0o^:�yr(�"J�H���(�	�5#�l_3�y�×4�(�Ԭ?~ԜT#C��y��F�(�4	Z�(�q��(�7���y"hE�y��xCb��=f�,m����(�y�j0V
r�z�iҚahH��燅��y"$\xW40�2)�<B�䁘G���y��	�0�2`*�
�h�C�C2�y�`;�69�7&�j�Z�rS���y��O7�b�Y���+`���Sd���y��ULYsw(U?_W�Ԩ��y��?Zq0
 ^�|u
!bW��y"H���5;�GCv�e��!�y�	�iOv�p�
A+O��C%G�y��R�\�v09]ن�q���x�6B�Ɏ_���+�A�-HJ���U��6h�C��+��xw-�%ab�򉈇=C�ɾO�L��L��_BnD�5)�\\@B�I�K}�|S1�N]{T@�ؿ"dC�	�-�M0��\46�,���F�RIDC�I$GON����0fRݛr��C�	�f#����M������é@�C�I�m�ԡ�f�05���Id)�V�C�I"m���RL�:<<��%*�B�ɩm��q�i);� HEȃ��RC䉹%�N��.C=w�X3�.�?U^�B��4S����>D���Jc��B�	�$@��j$�ާ
غy��$��cRjB�Ic=\pv!��l�rT�@�JB�)� ~Q�+W�k�ypc�1rd��@V"O~��/)-2Tcd�B�Z9���4"O �a��^���rB��!M���5"O��2�
�F�B�5/6���"OH=�G	�v䨜���ɯ[\��"O� �"X�	���R��
= ��v"O,LK�j�-��%PT���:��t"O�0HA�&(����?ZH"�"O0$3��	�N���qe��k�`�2"OH����%�ŋW�M�Fl���F"O,��eY���Nόq^���"On�cA�,t6p$*���f7�ظ"O�|����'_�> �Qq��HA"O�@ �F���TI,"�B���"O��R�d��SL��Ӥ� ��pP��"OLT�u�K�,��!q%��=F�
��W"O$X�!A�DKfqcԃ�1g���"OƝ���̯+}��PVBe�$8R�"O$�;V/X�(TNyR��hDA#"O|l�d/_�4zi�d�َ'�M��"O�4��Nޱ<p�1��<_�PŁS"O�!pҢ$�|٠'�\�_g���"O��!�'�{6��2a�L����"OB�8E �n�9�T N7Q�8�"O��ZRȟ&	�`8@�ϻ	º��"O�̀��F i��W��%̲�p�_m�<i��	��P��@Îp��e�Sg�<Q3�Q��NDz�"�^=$���@b�<�3��O�,U�,˂Xd��u�b�<��+�91�A�5��v7j�Y�H�]�<�d�_
@�b��`EZ�x�|,�� S�<�ÏM�!��gËc2:��$�	M�<A�o�	:����ÆI��z6KK�<�à� %�!c�� ~�&*��I�<Y��ߔ("��!�zf<��6��m�<�W�m8���3d A��l�<11 (�x�+ՠZ�\7�5��XA�<Y��#L �Y�aM0	��h#E
�|�<��޿vp�p��/�Jl����@�<����bd����R�V4u�z�<��Ȋ1�40�m�WRl�E�{�<��!�7N��kae�B�P��D�m�< f�4k����NB�*��+�s�<�����������Q�/�r�<�"^�z��� 	F5p��Avo�k�<�@��yW`�[���3(�ڱ�m�e�<��%@[��0��.�t��p���\^�<�uf[�V�PL��nN�Ce�kS^�<	�B�\� dK�1���'��[�<�V�̞T���Pm�"�h��pd�P�<��G'���8�J��v�
e�"Se�<�s��l<h���̣{XH��#�w�<aB@˂|w> y��� w3<�⁯Em�<�g�вFм�p'D rc:���I�p�<�Ϙ<*��"'k�0<��12a�Vj�<����>�R�C�FX�t���jIj�<�iΉZ`6�c֧N$8�)tL�<e�+c�f��4"�R���*�l�<�rlH�G�zt/�9S�	���i�<q�A��C����,����p�Rb�<��g��/���h���,�x��5B\�<y����d~rx����6{��D	Э�~�<����;G¶�!P�Tڪ���&�w�<!�&�LȠC��.p���g�_�<� rT dM� *��1Z������"O����N�p�,8w
�s�v���"O"hx����BsDqj檅�lr$��"O.99E�Q�"�`&j�~n�U"OlL���������׬F�)Pb�F�<A%�S99@�3�3� �9EDA�<��*"-^��`��rԻE�VD�<1�NF�[�������2�~@	�I�<�Ҝdf���L� �|�[�o�<Y�!����8 F��y;6���O�<qB�(��K��E�L�PX�kr�<I�e�"zSJ��N�w�8qQGPw�<	��E6&|��2%��H>R�����u�<9���m� y���F�a�+�v�<!��}@<P� �<B~pq��ퟰD{��	�%�z�q�-�h���0R�ߚ&�VC�Ir0�z5f΅N���x%)+I�JC�ɂ,� mB�U'L$V��&�t>C��R^���5�RI��N�~C�ɼs�D�bG�h?���)��B�I�H.�d�m�*.�:P���W� _�B�	�|	�����lKV�R�S�0�΢=���hO��A&�J�� I���y,A#i�O��tG��'9�5�U�T�\pS�Nd,<!��'��p�F��_�D�Is`�`m��:�'�H�!$*Y0Lk�躒"ˉbF���'E��C��g��uz���M���	�'�t��F�߿�$M�Ej]�Fz)��'��,s��ޮ{M����lC)<�z}!.O��=E��܎]Z�(f꒓<�@��,K6�y�(o�Y�G�O#��l�QE��y�^�{+v�q��N�0� GR�y��+�������dM"����yr��%P0;�+���M�?����Ӓm ������!�����2T���c�V���Þ9}$����̏'f�`&�0D{����(oZ"7���vĨ�$���y��e�4i�l�1P� �@ �yG�X��}���l����Ǡ���y�GR0 ��t�5���1�(���M�+�yrF>Dl��#�,T�'�A���,�S�O���k�I*g����0	�F���J�-���%�����s��!�ȓp���N��Z�s7�S��U��< �12�E�-��e��h��g1ؙ�ȓ6`�#�!�x=yd	S8 ��8���ҥG��hɚ�FmM1F(���ȓ��ES�
��D_2-S�1EU�P$�tE{�O���'�F,�d�+v�ا�ִ+BB�I Th����E�J�zx3������d+���3�V�l2<�����soF�s�e.D�l1e@�8��b@�3370�,D�89�	���tqx�-ˤ6� %�m'D�4���P��@1'H��,����7D�x�!l߼^�^ ���I����g4�D%��?Q�ON��v
J\z�-��
ع��	�"O�-i��2�^�&C��T9���F�'�!�N�7���`J�
X0��+U͋b!��ņl�Lj#H}���1��Z!K!��j z�A��Z+�,m��j��4`!�P�
јL�UF�J�>4z�*��gG!��7�"$���$� x�E��@!�Dʜ,�� ���bpv�j��Ɣn@ў��,��uP�˜$rh-+�i�� ̈́B�)� ���㍔����ǌ._w� W"O��SFL^�`#����@C1~hY`B"Om��(��G� �@-���2"O^�����)����D��>&��<��"O*h�@�4|�r�@P��)g^*�"O�hx���9/�ѱNE�R��|�)���4$nҢ�@cN�c�W>�h�*O���dh��+"��360�(��D�Zc�%D���K�"`6PHU��
A�
�J�!>D����!f֬���-z �r*D��`&�צGe��ńL ���'`'D�e!E�����w�l�Q�%D�|�4�\1@5b�k�
���� Q�84�L���b�4P3&�P�.ei���wy��'K���&��Y)��I�A�a��-!�B�N��!r�<M*�c	"�B䉫DӐ��3�6i��#	�nC�I�m�B�#���c�n�D#%hC�	-�� ��$ �z�!�&�2�ZC�IjB�HI���1.�j�I�\���ȓd���0h[}�|%�����e�~��?	
ӓd��󗦞�U�Lpj55x��ȓu7~X(%`�j#�J)N֐�ȓUw��c�JQV�x,��g��"��	�ȓ9����:UJ��q�\�-~����L<�7�	��D��&+4�ȓ2Z�]ӤZ�qQ�ݙa��E{��'�`QzUA�OB&����%�|�(Op���٠#V�I0fb�I �ٲ���!��;I��pe��D�궬��V!�DϷq�Dy��ʉ)p��t��1#�!�D�  �"�E�*U�i�eF�[�!���Id�!i��1v��m2q�/���Ο��?!���j۰�j��a�8�3gǁ	�?I-O~�O?USe@_V���[�,۬TʔP�taf�<�H�?מe�h�&s:,+S���&��F{J?��NSr�T�:b�s�F��k4D�d#�^�?���H�葾n��H�q�>D�� R.9{W��f�a���@ <D�P��+߈� ��@�C^(t�O�<��B�0�� 
d�0&���S,p�⟄�	L���芷j�PݡS�M�.��]���0D�d���Ѵ|�pLi�ʴRK0)+⬲<�+O���d�,d����T�\�C1v�J��_,<0!�AH�t�22a�9]1��ɶ�Q�7�!򤋹���A!c��o;��ar�Q��!��Y4w�|T��΂9-���0��)?=!��¾Tɶ��'B�!�u)��ǅ4!򤝶3��=����Y�
�㭐>"!��B7ah24�%��3�Hl����]r!���"e�*qL������Q�!��� hk�pY��f޼����Ģ`!��c-��`5��5r���x@ X�	!��W:4*9:�gެI����!�$\J�ʠ�bIsp��P��؉m���)�g_XZf���Z�K�ɉ<�͋�'Q���%bO�Q�����$�&�v���'xP:��Թ!��@6�:"~�9
�':"Yy�,�p�dMSuA���k	�'Q��g&AT���#�B�W�d��'�l�H�L�.g�ֱ3�f�;}l-"�'��ѵG�-�
��$w�)
�'�\��'픞B����7ț)t���'G���*� b�Fpa��F��L����� ���2
�@ǭf�$| �"OVԀr���:��<:6��"O2<Ȓ�.��*��W:c7ؤ@�"O�,1�aI<< j5��7� 5��%�S��M�6�4��@L�/}��4�v�K b��'{ў�>��Ƕu0��׀�a�ܽZƹ<����	WC�,�#B�*m��`č	�xZn�ȓh�Ԍi��@�B��R��4br��ȓ/�|hs�ƳA"XhFş1l|:=�ȓ��r��%*�(�gői���<ZȊVĀ�a�V�S���
�%�DG{����B�x�02GE�(sXHy����yb,7\��$����pV��B̗	��<�����	X|A��t`���&�Z<6�'6a|�(�� �~8x�l�3<�@�F��y�F�)!� �0�Ɇ�;��I�\��y�.�]�V@a���6G��S��Ƒ��O�#~:$l�,/���Rp��[Pu!��	m�	Y���O���'c�6I=�Jr���+R�l)�'e�P;��I���9��o��Afȓ��d�O0�4+A��>>f�����v�Qx�Ȃ|�IN�Hr��D�dU�&�A�^�	��=D�Dc�K3Y\T	!+�	O7LM�3C'D�䛁ψ� ,�I�3K�<���&����l���M����i���.�|�r"O4t�bƁ`c���-�#n�(rO��6�.���R��`ExQ�Ox�=щ�IY�FP�����F�cD�fv!�$��E�9�`�s��m�F�3_!��S#�4��/�J�ci�#\s!򄚊����� �I�t�Zchü"^!�D�pO���"KR7)�؉KW�V��!���T!��n�w��y�C�P�!�$�*8(� ��AQ�h��$��"2���f�'�ȭ��G�:-<�`F��e&� ���'�<Ћ�d��\��I6cbY��'�P�T��DZ:�`A�*T �'G<���D^�v�����?Qdy#�'�D0��I�`�D\Ȕ�F�3Q�4����hO?A�R,���Mj��' �@DyuY�<A0��%ZטY)U�U�Tצ�Ŭ\�<��Ǒ�����)|9���p�	e��"��
YЬ��%�R�yE�6D��8P��8��� NG#8����0D�LHfd��y�TS�G	k��X�&`<D�l��J��D��"r��z̄����9D��KD��;@}�X��d�r��`;D��t�^�Fi���6|��.D�+�+��l�̲� ˊXbM��B8D�XS�[Dz&�j#�O[N��ҭ;D�к7��&$��\���I<l0;D�ȃ�#D�=����,wjL�`&�7D��+"T.t���!x0`X�`:D�<�b��"��-y�Μ�'����g�9D��P��*�Z%�M�r�x�H�`9D�L�6�	 l�8�gBF��`��Q*Ox����Z�J��e!�r�P"OJ���`���-�ح��N
�"!�®����ȯ,�@���΍�`!�W;�,���`_� ȸ@q��Ӕ3�!�Dǻq���f�����$��X�!�D�^��|�d'�%-:�|3�a�M�!��0*���H�7"@f�˅GW!���',�I	� 5uR� �Ìڷ B!�� 8\��\@�Qq��I<D��!�*O�%#G�]&@-N�qՇC�C��U:	�'����� Fd�ճ7N��U*O������7�*3曨
� i�2K[�B!�d��]AX(z%���F�,�� �!�dČs�Г1��!|��[�	�E�!�dM�8��	Ёì+�@(�5FA�@�!�D /C��5Q����o�j�3�
3c=!��'-��hV�Ǻ�D��.3X!򤑛�~ �����X�>�z�,�0�!�S q�9�u�ߩi�zx��(Y�!���֠�a�h]�#���`K
E!��9D&1XF�����jA% �	�O���$ثu�hr�-*�*����~!򤅊VAT]sfg
�b���Ǝ�
!�$�� r��@#�M�@(�df� ~��'�ў�>u���v���H��u�vh�=D��+�Z"�\�3n��k\R����:D��Pd��	T�ЅӆHN�Z�x'�:D�0������I0�9�"�fH ړ�0<-�2j���P׶ �A�L FB�I�P�=�2��r�{�ύ1f C�ɵZ&hsQ@	'눥�ӂ9P���F{J?� 2�'8�Ұ���X���d1�� D�<��I�kM의1.Q+92�ܨ�j;D���LD��,1��έh�hU��e;��0|�T` /d���S�Z)�$:��]�<�2�N;J�����H��~̙Kn�m�<ღY2Q�������H7���"_�<i��������)"��z0m�Wy��'��OQ>)"���V�@#�ƭb14M+q�&D�\��O� /���Swl���aª/D���T�W>���z$䓧~����w) �	Y����>���Ua�I�f!��b�4$�˓�0?i�iS�ctz����©�����o�<��Ú
F3$p(G�pE`�����V�<Q���G+B��ĭ� d[4bEg�<!P��1Jb����I�e��M���b�<���>�0��V*ѨF�����\�<�gO��o̖�)��_f����JX[�<��i �%@$$YVGQ+S�R���k�	H�H15IB!v,��`��4'�M�D!5D��{E*��x��%���1�4o74�p�Zy�<36&F�l����V�!���(JQ)�G ~slq ��TJ�!���|^6�x�ɏwZ�m��ˊ�F�!�D� N�qA���K��X�7k��=�!���c�Ԁ��X�P����IV
�!�D��x�8,i�PB
̀k�'>8L:�Y�.# U�6��5�ބ�'����"����0`���}9^	�'��{�p�"��~�"�cU��+>�>Lє�.D�8Bd�_<Uh� ˍ`�b�X��.D�,3rfX=	�:��!͝4:�F��&b1����?�&��Ș��8:��&dn����_�'D Pq�ݽ	uZ����5gD�;�'��T�%�ژB@���hʢ~�V�"
�'2b����T����G�]�?6h���'�
8�aЃ%��(K�6�l!y�'��:7�ևԨ�;�b�4��8�'JX��Fπ�2���ꀼ��@���$?Oz�����.��$	=V�`�R�'��HJ�"w�8�Òo��#�`���/>D��HG��;7�z'%1G�p��6D�� �0EO�hހZ�`�5�}P��|��$�O�b���Ҍ'+ܜ�QL�,"48U�0D��8�)�-�R��j�:Nԅ��/D����Ї^��pm��XL��.D�<�S
F�~�p]c�,� ;������&��0|�w��F�J]p��̂('nh14&^�<�Nڮ3��uU��Xc����KV�<)���t�J�Kg�?�����(SX��0=i��=^�5 �ߎ!�hd�7dp�<	P��I�f�[��G��-����p�<y�*�<!O⑨��� �����D�IA�S�O�R�3�	%uZI�UFU�� ���'&ў�D�D��`�t	�B #�.�S�"C3�y����5B�0CanP�*n� �ҷ�yR�� 4���%�?)��4���ľ��'�az"d�(D̣f�ٗL��@e"؂�y�e�Wa"�����v���b�y���~���ѲiX ~��q��M�%�y�K�aN����@�l�<E ���yrB�5���	����d6��@`F�y2�ω���j'W+(��wα�y�e��5Ҩ�J,�7�9k���'�azR��*c�Q�D�5Cʪ����.�yB`�V�|���O�#7 ,�VD^"�yr㘑]"@�v�ҍ=�֥��NS�y�ڿ=TU��&:��@&����'�az���~�SX;:A�,,�y���L�Դ�C�I�6(� �DD��y�&ϻ($�HB,H�2�8�(�� �䓩?�� � ����/&~��=F1����usT�h5eQKOh$QsA	=�\4�ȓ814i3)j�l���kَ��V��AD@�7Ը �4KԾX��ȓ%�.���^�+^���$j�9:t���ȓNT:A!1l��fl ��8T��ȓ �l;�b2Kb�7�T�p�jy�ȓ
2��Ya��dN�0��(J����38\!p��yFb�B���!Sx ��ya��ҕ�$�Ƒ
�α?\���	f~B��]ֲ�(f	�H�~5ۦ���yöun@�ÆϞA<��{�MN�y�`M
 g�UQ�38
������y2J@5�hB�l��<��K@��y��*r(!f�>I�a*�	O�y�˯K,�}8�-;=�ΝJB� �yrbZ�%�@ȕ��5�&�rB
8�y��I�J�� �c�(����H��yR���DL�0fƴM7�#����y�+�p;HU����>x�SC#�y��3ά��!�6)�$49A���hO��ĝ�	7^�y�G6��s6�Lq!�D�L�
	GhX#n �˥�� Gp!�$L ���'S2e�lȡXy��"OP��s��E ���ڲ`t���""Oh]�GC�;\j,xפDk��[0"O@��k��>�H��͐)�F�	�"O� H���KŠ2��e� �'��'��)�'aM�}�&�AB�U�䡃�v<��'�J��жLW�11dH��'���*��@�j5��Pj^�i��'m�u)$f�M���aq��Mo&]�	�'4����g�=_.��Ȁ =jB�y	�'�&QY�.9~���Z�F�n3	�'3p��#��,&�b��@�ǆ=�0}�	��� ڝ���ܫP��RV��t�Bț�"OR��7�͹G����LK�w&�}	"O�H��D�7XB��KI_66$k�"O���C�;I�����	�h0��$"O���`�2'r�"�nF97(bh�`"O��`Z�jk@)Aȇ�G"��z�"ON�Sk�%p(i���{\�I%"O�j4�&?C,eТ�-0�"O���5FJ��P�f '>��@�"On��E�D��B�E��)�"q��'���@ܬp2(��E0	f�)AP��<��n -AC��i���xU����؄ȓW�z��!(|=��Pn�(��*�r���b��%(,���	=]�E��v�6 ���>]lDXڰ�X-XTy�ȓA*�[sT�Fe��ZE�AI/<�ȓP��r�H�O������	t�d�ȓq=�}qn�(T�0��S
�N ��9=��J�Fڈ[ԍ���^�u��M��]�5�:>��T��;O-(���%;��s�
?&�'P=q�bd�ȓI�}���#���5 �"4�����rq]����y�h��bs`��ȓ��9r�&σ}��h��e�:8G��ȓ1|��w[���ڵ@��mG{B�'W?�;I
|��tB��F���b�:D�H��Z.�!�VBG*;�m�e�=D��b����HzF����y@@�l1D�p�1HYcl�A�d�*h���Ua�O����OB��*X� �BĻYw&����֚;�!�D�=:H��-���CcnK.�!��������^�g�ԁ`P.^�q��I�`�?E�DN&T��	9��D��� �'u�<���ο.dz��Έ:�)P,]v�<���H}â]:U��P>hEY�'�sy��I�\�<9 �G�n��l
��)Z��# 矨�'+�y?O��$�'nL�9��ǱWAR<i�"O�`���I>��t�  y X͂6"O�M���A�F�paIY�[��@�p�'��@�)�''[fi+t�?/k�$�SC�@e0�Y�',�1���D�
�x�U疶6`��
�'_q:a6jX�ԣ��.���
�̘'28���(^fC�3� �"&|���)O��1�O�@h��ޤE�j��&�=_<A��	D�d��&��^yh��'���FhH(Q��3D��Z'�J���\{ΐ?����B4D��sW�S	<��)j���+�ɩl3D��p�났?��)�#	�l@���G�,D��(��W���)�#��.��i�`g(D�`┬Βf@�t�� �9\����2D�����vVAƣHR`�5�BB2�%�S�'LV�5�sbF,x^�exs�N�x
�`��`�x�´�Јu�}`� ݥ[��$�	s�'Y?�1���	5'�3gÜ�L�8�G$D�t[����4
����"D��{A��mr�!�WN�3J3�Q�g"<O#<y��D�~|"҄:#��!R�C�<au�3=�ČY�C�2R��j�g�V��hO�8
Ѓ�\�*t��㰅%'����qm�b�E�0	��<+�d�; �����A�|�ړ$R�Q��e�ӏMp(M�ȓH�b�"wA�0�� �Eوr� ��U�F��t	C�(�[��< �uF��'>�Фe��R�����͓$!�=q�L2D�� >����G�$ReXa����:����O<��I��^���	�}���6��Z!�D�	M�.)p����Ƽ�����3Y!�Ċ?p�yI�	�+�&� n�!���Ib���4�X��{r��,�!�dW�"���1U�j�b�� H!��C�{1Hh2�\�6��K�*/4!��%Mrm��љ?9��0�.,!�ZhsP8���̝?ؘ�5�8@ !�D��kp`��r��[P�kC�-n!�DK�{T0�EE5C��Z���o!�ۜ'��ɚ'�.�0���O\!�D�o"�S�Ƀ*.{���.J�b�!�dž[=ލ�pMю\[�)#�m �&!�J$�T]�DҚOA�2�Jښtџ����C~�O��+�S�!�� ;�+�R����'/�tHÂ�w�P��U�?J$MP/O�O�����v��=i�ɜ&0l��@��!��#����f)�+j�A�Sf�r�!�$F�>���v���ayi#�T(�!��_P�-��=-V�Q����!���
N���٤iU�i��D��"�} !��=�(�Ҧ��	|@9xA��!�$&#A&!@�数qh�0 ���T�!�dH%+t��b5)T?RgR�A�I�!�d�ek��'�n-��R�g9O�!��%PY�)�R邳���'48!�D�����S'.�\�Τ��?2!��M}4��u@H��̛���!�$��r���)v�V0��t�!�Dۑ,���v�ԹJ���HX({!�d�q�x񳴧��<H
�j�׍6 !��p)QT䍬8;���g�PF!�U,ZG ]+���"L���1>G!�D�)_��[�%o

Tj4$�)!���&�h�%���EC�6w#!�dG�.j�Y(��Ԓ�������{B�G�/]���ê�=/X�J����J�!��)q\��`I Ha{��<\�!��W0
xP���T9P��5�ǃ;w!��_g��i��ڈ���Z'��6k\!�P�n��Ea�)�=
�	���Q!�䂙)��L��A.s�0�5�3UF!�Ȅ%��d���[�C�>J�F\�7!�$R�$�@���Lc�t�&��k�!��B
}�x$�&dZI��A�M)"�!�Ы?����J�G��H�b��D�!��M're꣥�N�hf
C�<�!�$A3=Zb��啍%�L�Q�'+}��)�'-`ӀA;K�$d�4�]���	�'��%��@�x�B�êYg!(�a	�'�r`a���i�X��*Ěr̚��'Zl����19�ЉQ$3s7b�R
�'��PYT�O�G�\;�O��;qެ(�'�����*X<�p)���9@H|��'����e�_$uY���O$I�n�����hO?�: h&&P�y�����[?~M:�Rk�<Ԇ^��<�c�`�#�	��
L�<iP�#dݚ�C��> �eaC�XJ�<�g�".����U��{�0����~�<��P�Q�`�LқFvD!2��|�<a���r8J�	*�"N��3��m�<	 Nd�`�Btf��,���{r�jx���'�d����Q�\����`�C��x9��� �Y�
-7Œ��"��TX�"O"�z�Ê�-��nR����"O����f��U)!n�̦�@"OB�� ��x�ę!�=�b"O��0�˄4��<���5R��<��"O��q�M23����/ؖ?�.�Ha"Oz�sɑ�k�f�'��g5��w"O<[ԓ:�l[���t��"O� ��KR%o)8�{��[kV\��"O�iqG���x֩)��[l9
E"O� �E��	H�u���V� C�Q"O6)����3�� ��dߕd�(t"O�P0�?N&@bd�����U"OdhA��%�r� V#�.���"O(�H��9=�N�����'Mr�8�"O��@#ǂ$�>=Q��i�"O%�c����ש�y �,�7"OR��&*`�,e��钺_�d�r"OlPS%�4l9b�腨�[y�<k6"O,ZG��(62��f�7ql��"O��i�+��͙r@��
r�D3t�'�!�� P�#ߌ�.�!P%���!�_�<�8��ŕ�r����S$!�W#`��Z�kJjA���Ƌ�/!!�*5F9��HU ~'b8y��/ !�PUl����+P��xB���\!��/aW�q ��C(#��-�!�$ŧgQ�dW%@Y���g�'y!�d�2H�D;��=x<!��e �`!�Z`����No΁�7��B�!�-KDB��B4e�lXJ��	�!�d*mH@��ƅ�"�xk�Iػ5!���n��]f���-`�J [�!�䑑-BP�A�-�D�Ca�ȓL!�d�5��Y�W�� :�j4c0ɘ�VU!��J6�8�Q0�YZV��GR� G!��*���ք�E��&��K3!��=�xq8����m�X��CőC-!��3J�6�5�.z�P522�Y�!����˵M��E�\X�F"ۖ9�!� �&L[�*��+���2���B�!�$Zn�� ���riZ]��˝��!�
_���X������!�!��ܳ(��ab)Z<W�58��Q)]�!����i�C��uX�e�<s!��[���3��׷ d�R�#łD!򤝛^UiL�&k�%�$"�#B!�DԆn�"��KV�:0˶e�0,�O6��Ӎb<pa��BtHe����8O|!�.]ep��^{�ݡ� �(I!��@t��� -�C����	�� >!�d	�E�.��Ađ gX}�D�9#!�@�e�����rZѻ1���r!�d�||d���%��`J82���q�!��aC��"qj��{?r�ʃha!��Ь]�r��X �Zt@ �rT!��T�B�V`p�N܄��x�P �"s!��a�IZf�ۿU�ѩ���2^n!�䎂f����\�0=�L��-�s�!�d�;ШT(Q�Z�̰
��p!�ă�9��ĺ�(ʅL���Kd*Ǭh#!�đ�J��|`'`�~���1��UB!��5HM�5�D��4\R��P*�!�D�2�|�1D�_-���Ӡ���!�� �q��G�$�^�⏛��FT�"O��tc��{���� ˹Ix���f"O>���Õ�0R�Y2�R7nB%q"O�X�a��� �V%~�1f"O����/a�0J�͓ x�xi�"O�Xd�߽o�V�y���ĈAxP"O�R�o^g��r��L�l��"O~�g��&B�u��ƒN� ,�E"O�x��j>A�6��d�?e�,ҡ"O������m�р���`=��"O�xE�N/��� �.Ӻ�[�"O�U�#��}?t���Ɍ;�P���"O|`aY9�����HS�,xe"O��8�!ڜXQ���\���jq"O^��Q?R��(qC�)@���"O�M�eMP�g���,�+�H��"O���� �z����R���b��("D"OH9���L-Lv�I+hS,r�r�"OJ�� -W0U� �'O[{��:�*O�<�AA������ڸI���(�' �4�1��.{
�AFe\+��Ց�'t�<B� �~:��f��%�}��'�b��'6��$as�� ���q�'��M ���_� <��@�TP���'�Ri2/��8V�*vLO]�.�c�'6���
�K�0�� iE����'m�aa!��?)n��m).�2Y	�'����J�d�LeZuǾry��'jB��!�a`d<�S���i���
�'G<UkA�'t9Q���e�pu��'LZ���o��^Xt��!�W�$��'9T�c�O�S8�;$"�z:Ĉ��'nyc�`(
�Bs�Yp���A�'�LdC�O>4�D|y��f����'ƕ���B�	����Dȉ�Y�x��'�-``�I�@���ÇU0O�����'�(���.[�Y�ŅFv@��	�'�@���E�o�b�p2�ܧ:�xQ	�'p�q��#Z�,��x%�7fv6��	�'�.����^�����@,��s	�'4��!��<:d�� l��1�e	�'=@�J��C&�D�a�I� C6ƍ"�'��!��'yĨ��nV�:�\X�
�'�&���g�*l�'�*+E��	�'|���?S�V5jb�˗"�Ri�	�'Y����t�q�*Xjl<�`KXN�<!�Kΰ9r��nN�dL�u�N�F�<1��5Z�L�)��0�VLs��NA�<�Å�$:�by�2��CB4]Pa�z�<!"�R���x���^$@Qx�t�<���79n��y�(��CY8}��JSq�<�FZK�<�s�JO(^���k��q�<�tI�?OHZ���h�V��l�<A%A�$�D��eb�6K	�Z2/P�<�B_4t����n�^�yrIr�<��ĩV:�0��E�h�j���j�<)�F�PJ����҈{�nL���f�<I�a^�[qh��S�s�M(TlWx�<�R��3��eX��/-&0H�lJ�<QS�2"����Ņ��h��"I�<a`��W�!��J۰b����E�{�<����n�D�2��0��l;d�z�<9�]�,2�hRg̨L���JG[�<�v!7
��#�J*&$բ��Pn�<� 4������(l��f旳0PN� "Ov���nRl
����_�R&���"O�;SC�B�]���� �LS�"OBH��j��^&0{��n�$1r"O*�㧯.Q�ɨ4�ŵ.Қ�81"O�Qs�$G�.�|�R$�%X����bǤ�E#ԓ|i�p��(g����E�Y�&����&4��l�ȓ\���,	-h0�P�ύ!B��ȓ<u�a����qT�1PqZх�2:�5��pl0�W���7�����y@��ᓅ�(8i�UZ��	� ��eJ�i��+�nG�Rv�^�g�Ňȓz�\hقCD�o��5�ـM,b|�ȓK�F�Ĉ�ۂw�ʿ�@�ȓo�ЙPOI&�����^9`���ȓC+4AE��Kw<eHݳ�>�ȓ%T
��*U�K�|��dQ6;�x�ȓ^����sBA5�~�k�ˊ�u{ԅȓ3M���1��RA6���$�#�Hh�ȓ.�>����e��9�(ʼ���g�,�T&S�숑"�1A�T���_�"L(�����-)lC^ڐ��ȓb�t�sI�5J�dՐ�.C]�ȓ|��q�g�fa7d�)��\��n�@�<��GC�0� �!I�e���(7F�S�<Yר�z�t�a�N<pbO�j�<����=$Զ�فI�;d`��Ac�<Q OШ.Ʈ\Ö�'���� �[�<�o�N����eW4XC�/�N�<�	��bt�� 7��>7tބs1�\I�<)��K�a���d�$�b4k `F�<�1J�B:��TK�A��T��	@�<�pOԄ��lz6�	`������|�<�.֜G��h�l^ ��xxv�y�<��nY�¶����Ϳl�N���i�r�<�@��A�`!��!�����\p�<)�B��CT|p�0	_�� q��m�<�����`�R�FD�M�0��_�<�@$ÁvXeu��r��Z��Z�<铨<Q��B�-ȃ �0��"a\^�<��$�=�p�ɐ̑�p삽�QS]�<�(	�?"Ġ��M� 2<��Da�\�<ɖ�ۥf; �#`D�n�^XQD�q�<`��7W^�()��T�l�
Y�1FAo�<)��BkV�9��M!BWq@%�^_�<!#�ξB�fh�gȋ�Ƃ��X�<9g���C�|1yA�L����S�<�	L�o����@)�[�����*�i�<aa�jd�l�Fngqn%c�Xa�<�c��7�H]�!'�*lL�H�.�U�<a�@��{%ب�w�(�8�3�F�<�b �Y��t��@(wJ�p)2�M�<��FYC
��ا^�0���b�<�!ND2B��պ�aW
-����Ɨu�<�Bg��!��z&,��x��l�<a��Ӛx^� ���tj�XfbJ�<���9M�-(��܁tΘ�@�I\@�<��	�=W����WF�DT4��Fz�<�f�qX��P iL
9�4�l�u�<�R<+��r��f��t��aIj�<�c
�
}�5d.ڏm�f"!hI��<��g+��+g�Pu��0��مȓ^�P5��0m:R� �)@0SI2q��S�? �љ��2]h����n��˳"O`<���S�X<���"��!ct"O��p��!��q��C�-�"O"8�dk |o`˂L�&Bġ"Od]1��ZbH��*��tn����"O(l�W��L���P)\xP��w"OP�j%,�N�0��'2jy��"O&���Lp��q���4���"O��`�f�$�j��ƍ�,��)3�"OdQa���)�T W��0�.]��"O��Ȅh�5q��=ׁG:B�0\{�"O��Qt� ":&�u!G�4�N�"Ob�hEz2|��Ƣ�F��i�U"O6ᒂ$_�	��p�g���/����"O ��G�w+4�9!k�8B�X��"O<���W�H9H$�%�[s�3�"O�ha��A�1(�QR(��4��"OH!Q� �	Up��gF�<%V�UCt"Of�뢈�2��y%	wF���"O�`͒*H�I�W��6?|t�#"O�@xs��h�BP� ����"O�ahi���M�6�i�2��a"O��ؖ��m��#�c���s$"O�L:ؘ9N���#��|�1#��!D���p	�v��A�C�#��]��',D�ru*x� �L30Z�mz �)D�H;�D��1��HڦL�~���	�()D�L#���8r7�Is ���%�(D���v��20�a��#�hr�)�5�#D�Ԉ��J>\�JtB��et65k��#D�px�DA1jC������1Fb���"D�D��a!�ى�hP�R����$D�$�G��s�d|�@<#OH0��� D�$������V��֡��z�,���?D��7iP�g���I���"t1D����d��W���Q���Zԉ:��"D�,�`͛�&u��Ibc��!��`�v&?D��@#���*G�-c5�.Q�`��j)D�t�a�m	:yXw��[�� �F�&D���� �x4,03��P�QUڹ�&�7D�t���<.�\�uH��:R�<I��"D��1(D�{�x"���)u�T09�d%D��`d��cN,%A * +ьd�1�$D��Z�j��Y$0MH��	DFx�%�"D��j��p9��ZGDωkIb@Q�?D������Pn�](:(Y0�!D�К��"�Tٳ�jɫ:��Q��>D�@!�)>����F�7��<D���uCZ?~+z�k���Q���i�e5D��Ԅ���t{ �'Mw�U� (4D�ܱ�[�_��Q�#��R����E0�C�ɞ;و�2�F���fȒfs�B�	)��}y!@RQ����э�=N�C䉚V��|a%H��p���CdN�3�OP���B�U��Y!�g�UG\�0�FS)�!��2?	j����WNn��T�HNQ!�$�F,pö��8oJ�`���C3!�Q�S�*�Z��Jm�Ux�P�~�' T}��	%�^IA�Z5P@���
��z����v�dX��4r$@a�@��b�A��1D��{�`à�4��pA�#���k,}�U�<�O�"<A�l�/ �e9�ܮ"Fn�yB�V�<�6'͡ts����!�.C����5%j�<��f�B�V��H�Y��2�$�O�'-Bi�V�π 2�� ��@�"X�I;d}ڣ"O��R.�_�Dk��å	v$�ē>�'{�O�|P���K� }���C��V�"w"O.�Ht�R�G�vi��Q>!v�*��d���0=�a�T-s�:��Q��6"6+A�y/B O�1��)�.%:�������~2�)�'S��!t
�jŰ�8r��<b��?QM<�Ba?��4^��*� ��;��[bD͔p*�C��&4�z�8����Ʃ˜.��=�Óx4�y�5`ŔZp�9k撼na�����D���`_��T�M�8�B �>�#�!<OTH��M�7
L[t�՛o�n�kF�'ў��$_�%�H9z�-O�">p{�f/D���	�2	#����Δi%XaC )?������'�i%-� ��)����*@((�'r6 ���0w��яX,Ib
�'�,���(��kI�4Fj.A�'i
�4�ܮ/"f���e��>-4Ũ�B�)�t ˀ=�,��ud�Vⲽ���)�y�'��R{Ĝ*�*H�K�4%���hO���dK��xɖ�մX~`�A`�F6DP�W��(��Y9�'����19�EZ�bF�L��']!�DV!�(�h���%kHؽ� MV�d��'1����=��ڍWSLXS'@;W�D)��^o؞�=q�LJUÔ0ٰ�߄[D��H���g�<9d"R5y�4Pe�G$�X��Ha쓜hO�O ����F=I-2Л��O� Ȅ�;�'0h��O({BM耥ԎpL�u��dCV�4��ʲAI`c��ԯb՘!�c�$D��і��*Wf8B����`�أ�x����$�͟T����$�� ���BE�#E�7lO��y���=y&i�.�TIēr�'�m<h�}B�d��dղAڶ��5���%�NN��>�S��oQ���F�dl��#
%�)Fxr�)*�틋K	P�3��d.����Y[ܓ��'EQ���-]�xeb��^�U������n������[n�4Ц���]�xd�����c�e��I_}2���Je�W��Yq��� �7�yB��X�=�NF�`�Qp�L^�y��IP��g�8Y��r4�ȊE�����)CC��^��\����5"�����A��ʓR�IY���I��
ﾁ@G."}��EJ����#K�}b&�|}��Q-&���x�d+@q�N��y㈎Fj�a���V�0H{�f��?I�'�����W�w�r��2�|��	������+Ч�'�*=��<a��-:v�:D�|�7��$*����ް#MxlL+�	��$Er�O"���-���2�$��_��J�yb�)�S��)b����K�D��$OT	 �n��hO>�Bߦ\#�=�4*Ek}dE1#��<A���I�h9��W�`��YjdK�<�(O8���Vc��RK=[!&�+t�P�=�a|��|�k�:L��aH���5�@�q�^�O\�=�OPF��%.��(��#6����(d�'���#n�^H����ˊA쉡�'*���
�6$)P�ХP�)�{b����O6�t�R����2A�p	�`8O����v��o��b☙j��ǍGL$�l@�<b��E{��t&^���
�����0&υ�yrV�J3<��"��жt8� ����(�O�9�� L�`�"2���s�^EC"O�|2ƄsIU�EZ=��5��I��y���OT���`���fN�%����"O��xAO-[�y[�O�,X�Ľ��"O� @��aNդK�^�B9[}���c"O������ �\JC��_hR��#"O&���.�05�h������ک�Q"Oj)�7J�+k�� 8��L��6
��a�O%j�8�	W�#g��pi �(쳎yRK[���O��|����44��p��O�̵r	�'x��JB�H6�]����5>����w�)��<��J\I�H�e�P4���	%(�b��}؞,�0�^	4��вe�,wJ����F_�.-���	M?�PM^US2��R˺@1�8#�����hO1�:�O`��`��P����ϘYłL+4�	��]mZ}������[� ���o�iz���H�:�y&+��8�� ]�4�Ќݫ�����d�\"~����"%��2F�Zx����JG{�'�ay2��6�bEַ��Bb ���xB�U�PVa� q���q�H�{^���'x ���Q�&�hGɼ/�1jד5)tc�rUGԚ&�:�����zp�鈕�/D�,�G�lnX��R&�^کx�,�	Φ%Ex�x#6>�z��i|D{�c��'^#=%?�{��e��\�@���rX���n'D�� 0�G����#b��qo";wF"����'I�<�1D1|@�DpPb�P.�F'
w�<�W�#�D�� ��AR�£%�q�<��lϋUu��8�L	G(Ų��k�<�%��bER��ł?`�c��l�<1��8�vl��R;�;��Zh�<c-�yc�!p�È�I]`=���|�<I���$����7B�M��%{$z�	g���O�2$Ԏ��ېt��H�[9U��'"�ce��l0[��C�W�t��}�'�LR��@�ir�P�����J�ڵ��'{N)2�n�F������ʾQ�|�
�'7�	:��o���T��;r��J
Ó�hOfhXD�ˊ&���A@��Bx@�3"O,���϶b�1󕩉�*� j"O�{	��[����åSCk`�3�"O�[��k�Th��+y��%;`"O2,�tI j�j�թL1c}I�"O`(�D����t���Ά*Lr(0�"O�	��Ђeb�H�f�Z�\��"OR q#"�����G�I��h��"O��	�j�"|�J}���d��lA�"O�i�(M�>-1�J_�+Ԧ��"O����C]�3���*M	��PS#"O�]��-R�gЀJ%[N%��"O�<�"��Sٴ%{Vb�1.p�@"O�H�1b��D��q���J:ThH�U"O8̐�D�'E�\�����~���;�"O�"�5��̳g&�(��)R"O�3t�_�������G:�j�E"O���a�ӹo�1Ö�pĘ��"O�Ī�U�6\!�T!W?��Pr"O�A�SkZ���S���;���y��{P�DA.� �p�%)dy�ȓm9�=���KFJ<ٶ�Ay���ȓ��d��Z�v)揓<5Cm�����B��!}NT�7�<0C<�ȓ!�mPV[HTX��O m�v���Ir��E����u�F�@,�ȓ_�NmKdmK�0^��J���UwQ��Q ��RF��\d�f�γJVڬ�ȓ:^2	e��u�D���3��(�ȓ}6��DS1A)Ĥ��!��̇�S�? H�z4`��lR�pA�T8Y���A�"O:Y�	_/#�ʕ���+{Kp"O����>L~���<G(�@"Oq���:�����%Ψ�Z�q"O��	0@�"<�4t�c#�Z���k"O��c��3��h²H�6����`"O�-0� .����&]�>�D0��"O��I#�2�uph�
5I�g"O��a���MX�Ų��M
8����"O*�$��V����h��)�u��"OH�#�8���B�FE���0�"O��#�	�a
�D�Lt���"O���5%��V��}0�S-�E �"Oε{p�< ����	ӸN�~pQ"O��i���22���WiZ�%�y��"O� 7^�L�<���	�&$��"Ovِ��F�D1�d插F�>%
f"O��Mȸw J ��e�7u����'�N�9�/�,o��� ���N���re�+����'/Tt��D�s���`�'XԠ �'��d� E�F�Mb�'��!��'$2\;��
?y6B��"]ےa��'�~Eh����<��A8B�p�'���&��k��,�����ݮ���'�����ґK�&�����"��Y�'���Z�lZ�r|+�&�j�����'XT��F�ի ���Z�Z��'K4Y��<j���7쟉[��=��'�"DP�g���*��R�Hh��y�'�ҸSf��8֌p�Q7Q���	�'�\9������lx���S�\�@��'���{d��pr����`�=O�l�P�'^ ��Ö"a���'�*EMB���'>D@��K�7� �x��P�3�u �'D`���,��,i���S�*QA��'+T�jR�4"$P�%8 �����'ߘ�E���Y��u��?�P!��'U�T�0�[�0�I%Ɍ"A=10�'���J�^�l}
j�i�|�	�'&ZX�l�)��HHwaB�W ���'�؀ǄO��t�!4���'`���uA�,I~�`k�I�.�y�'���h��ϱ��!�tc���� 
�'�Lm�g)ڰ����T/̕i���(
�'���as���_N�Iy4��1)�n�h	�'�(ě���8s���V�@
#��Q*�'(0�R�)�z�2�i�����'�u���ox�T����as�'��ᣃ�n�L���N�:cV�d8�'<����eS=hr�b�!H�d&TQ�'��3��
�+�\Z�������
�'���5h�yB2�I��\�	Fm!
�'���!��/��" �?~?��'��)Qć]�t�8#�m*���'�4�CR X�R�y�m
�c�"���'����I��P�Bw��A8�:�'Y�J
�s�j��f@H�8a����'��L0�\��&�ތ*��a"�'3���=I�HA�����&?>;	��a%b�12%^O�:�q�HCg��� �� 
O@���2Ct-��m!�a�LQ�D�D]0Gp)�~�5(��{�,	�1Δ*`�Pe�AL�<��h+�ەe�$8�D������<���I1^^Q�#j$}��)�	�|�� hG�E����E�/(!�� �Lb�@�5?n�xeɕ�T������"��)9�"%�'_6-�p��q>a
Ԫ��왲	��B�r�J\�u;Bo,/������=1Enm��?�PYB�/w�XA3Ca����?�+N����b��(mb�>ыa��$t�+���1}d�]�@�9D���<�V���Q�*@�!0r�v���S/����"�>E�$ofg&ت�I��3��p�'�_��y"�B�R��]YV��-�lCwH����P�P8��&Z��p<yL�$ᓧ��}�Xa�c���t��8f�����PѴd��	���=;4�?)���&�*���A	xD3r�T� o��c�D��,��	(v)�nPeX��ϵDY!��Y�9�)ۅ��{iHt�$�1o6��2_�d$��&d1�O�zkL�Oju�q� �OcNջ� X�4�|�*E"OT�Su�̣{c8#1�M%3����>	f�\Jf����#���Hc��1��"��Pi��	��i`#�7YΔU[�'�$L�C��`�ڀ�ԏ�,F�@|J%&�%�-(ބ�O�lS�����ē��Z�gE���@����<��-�ēy�4�YuH�#��3'��F�L�Ӵ�S�P��\ �n9�O���h�+*��t 4E�Hj4`��'Vʹ���*�ܔ'D:� A=i�4��ď�+Iإ 	�'Ȧk��7#��ź��=)�h�CL<�%��9|]0���H9��^�)a��J,HT0�Eeǉr<� ��FL8a
�ݟ_������`5�qddS���	1�~؃��L<���9���Y�	��vQ =��ZH<]�J��S0���aK�GЈ�d٭B�$-{@�<�O��X��X�H3�,[ďI�_���'�l(	v�8��9j�i<�᥊X� �f�r�� :��sr D��DPҽpQ��P$~��' ��M�\��e�N@֔�Ё�:��O�bT��Ą8a�H1B��R"%������i�f\�p�J�e�L���`φ_J��Aa�g���I�l�k	�t�х��J�AV�*�3�ĉ�K�n�b��=<\�D�#� T)��X�6kȕy����|���%L�t�b��!�J͂5���K�E�d�7/�<����.[����| �Q���ӳm̘�q3`$t��R%��q[����>5���ٙ7�]ay���r�K56t\�2���+�H���BhH<1үٚ�$pi�g
�"�h�pD��sMz��a�
#C�;���-H��'��X7\�zt�̹+&.J�(P�;�~�B�Nx����*&D
��Ԁ>/���m'ٶ���"C�v�X�Ӓ>���I�M���
�L�=T	�ið'K�>�>������<�{��>�Ӡ
�<]#�J.��s��s� ˓6.&�pv��4_R���䗨^4�3�a��e�N� ���]�$�!L��G���)��K�J1��*�+�(i(���!A	�� @�	:.&���'��i����	W*$@k���" �U�J�@���\QOP̋$�3O[�m�j%�4���(4�+tu@�c+<���J�'�V��#C	! @��`�窩p�*Ҿ{CʴB@BB�RP�P��J�S�O,Bha�I֟G�&��С�!�x쩌�d��N��(�!%�S?-cX 86�ޞ`T�=y��=A�C�I�N����7B��i�@��3�˱Y��ʓ	����.�)ʧ?��N��8�)Fj\9f��i��?� YQbM�h���)�^6l�Q��<'zzӇ	n�h�0-ѫW�8���C�R"���dmP�1C>"֑!$j� #X|�Q�V��Hg�O����3N�2-��j��ѡ2$�-;��.lO�0&ļgP�I�7#�)s�́V>�@��f�"? hs�O0S���I,bݘ�+u鐋mnҐZ�$�X �*��ɼS���%��Rp�V�oM�d��74nF1q�L�?���d���<R�J� �f
!�$K�{�"��kW&"Ԍ9�G_�|��=�|qBm�{�1p��ź�`���X;�OdͻW�Lx��4r�(Q�	74�ل�I�/�m{sЌV��KM3�Z݁ !�2$W�4��A@����i�,<S��o
<Q���B#=9ǁܙ$�����b�D� �@��ah�Q���0M�����Ƶj��*�N4\�Q ��3kX6uzրR�-�(!3�������@	,���C�<-����*�DL��XT@;/9���ɱ|��ր�*3-��{��`#�̞*.]9������D�̞b��a���U�cVB��7� ��Fpƶ��D�!�= �
8n�	i�̛��TLY��� 6�$����Ywμ��� ��N2� d93����y�5�歐�T,��Z��'� BX�p�n1o�M5^���"����2�@�(k\d��պz+.�)Y)����&��M7T���4A41#s%Ё]T��I�BW�d*�jĎ%0n�
p�\�>],�	��B�H3O���S�ÆG_�t:�O1j�" 	\�<Y$T0D�?�ժBmɻ*[t9!	�3fpM��,(В�o�.f&(�HV#̯*%v�G|b�^Ѽ���ϐ�F�(�Ԏ�Iĺ��e-�K�]B䎀�L�>\�4�ˏ\Զ���P%E��S$a^d��w�F�K|�@BD��g��qj�O�x=z���'H@X��_��v��� a��80��G�%��|S4��:S{� OB�|pi���7E�����4U��C��<6��V�ʡ�EM5�d�x7��+�HOZy���ũ\�����'3T��S���?�2�옫rL���c��;y"��DM?˂����>��#�*~D���'��x0d���A�?O�0ق�� 1V����C1�,xYR�iYz�@�F�>^|Jy��.O`�I�E˺�"�U�QP�J�_h�p�5�U�W� ��Qb�W � �N�9YLXM�'� ���u������	v`d�	��P'a���RK�;=�$�Ig��SN
aJ�K�<,�v��#K��skr�A��f����"�����G\���S!v�L�#n9W��HU�92� 
�s�&	kP*��%v�5˰B�cu�9q ��>�N��o^�	#:�6���l�q�3o��$���

��A7$�ئ��'R��0��v���HH�4mk�-p�'���OD
=N�nڔJ� ]Smޱ�੠6���N)B��".�>~|z���,hD|؋Tb�*�F}	�$f
6Ċ.O��;��D���!��'ծ|둪�3M�<%���>W͚�h�4o?X�C��&&3\7�2% Bi�RM�w�0��dG)#�JRbT6.�j����	h\Ez!��v:y�e/�o�ޝ�'�(|�P�� yޑ� �rK�Z z	�c/3|<�,G]�/�\���bW9�-ˇ�#Uz�1���Ś_*h�s�2~>��	}�}�FÌ�{u�)�\���[��&�O�%�P��f��9@Ў'mN 
WHT=b_Ass'�,�X�� p�@�ƅ�45r�d�P�#gZ(J7����+,O�,�VE��}�+��GL�mXqDG7��=q�d^@zl��Gi�V�k�Ր"�*1��G.@~"Rh�>G�Vib��!htP�BD!Ǡ#�T�?���K�vN���$
h(} ��W`�'p�"�MÖ7�%�L�� ��E�.`Y�L��Ip �q�	�n��Je��S�쥋�'`���V�NUO�m�+ʾD�����H9ow��X�'P�)�%D'4M�Q�3gǫ%�2馟'��3J�n�cc�G����6Ұ�y��śjl�X��M�7�`�2�,� N	T����I���XSm�����Y��x��'w�����Ξ_,�-�E+D���Ԍ�e�h�̯$U���fӘ�X�Q?Pj�ѥB$���d��	�&��r-Z�on.�)≞,9�{�Ƃ#������M�ȭ�2煅13vA7��Q�985��JH<�V-�^��9�ɚ��*�eU]�'XR��fMw!才Q�Oa~�I�b�y�T5�u���S���;�'t��BC��)¶yP�jE�T��1s��4u��2L;�)�'4D��a������Y�EP O��1
�'�N8����=������r�n�{	�'4(�؄�є��\ՁZ�fPh���',KňWL�t�Z�nאhPT ��'hH8�tB޹!dy��VS�:���'�P�W�ݚ��y��a�$���X�'����6!u4Ekg�����(:�'\P`Y��&AL:@��(ӏh�
�'뎉 �R���zt�ڥF.�8�'����兤J��Hc";d0�3�'�n��OM�E�l3B��=yY�'*������e�	t\�����y��5=vh������(��ቌ�y�Ɗ�}I��� a8�� H)�y�ϏV.��e`@	{���X�͝��y��S� E2OƁpp��EC��yR.[:�,d#�M��r��})�]%�y"�>w0ܢ��B�v��[
��y�m�6d��I򱡅)�a�K��yI�<������)�����`�y�G*~,A3jל/j����3�y�I��%�i�A�RcZ��dԕ�y����޵��/_�H#��zT��y�H�
=���Ca)�
@�+�y�2n�^���l��8�qQ�@�y� V-`��-�#�[7('HH��"E�yR�M�V�h��4L�)}��3�ϋ$�y�%�:_4@e�`�-~Bqpt�
�y�� �V�CCU����t��y
� }�ň��rE��G�)��Q"O A`���X�!`�@�T��T"OR0�A�ܶ �zD� �>)��(��"O��c������ToČ``m��"O��������)b�Β?��eKG"O������$���Ć�� q6"O�9	Ԥ�6�^ ���P�i��R�"O~�x��е	�fP��ՐUG"�"OL��2'Q�b�n���k pԳ�"O��jRo�rXF��EE�\ ����"O���4���zd�3	��LN� k�"O:ɷ���u����&���"O�����U:?S�Pt�[����:�"OXDbe+@�$lh�׬^)TXN���"O�$��-��p �"�U�Y3``�"O���^�;<d�aM�I�+e"O�MZ���c��$B`틐8�X[�"O\�{v,[�*�b�&J,8�&�0B"O�-�����~O�����B���"O�i�E�,�4DX�ē�b���C"O�� �+��`��b�B�*:5ra"O�=+��F�.L�k�e��"O6yע��Lejq�U� ����"Ot�
Vb�$8v���	�r�8W"OĠ�0�O�Yf�X�A���Q"Od����Ar�сU�P�S�M��"O�ɴ$O 6y�ё ���.�  �"O�)G:bg�A&�6lrdXq"O$��N��sI�MY��X�{X9��"O��Z�"����Ce�4W1��r"ONóbʟqG�y��~�<���"O*�92��:n�!c��X�&�Jv"O�̙�%�J�ԙԇF�@8�%�f"O;R�N�(�b���MP�A�-�1"O�ܘv+��r��) �!E�A�*ձQ"OD`#����L�1� e�����"O(̸4�W�f��S�A!{��<�`"O�HB�}B0���3z��0r�"O���ܛr�r�'���,�( �"O�X).�4B����)	���q"O��� )Q�'�J�TA�8X��"O�\Hq�p�`�����C)z|rf"O:Q�p�2
���4��K=\`[�"Om��h�1H��T��9^+$ K�"O���w)_&	�  �,K�a��"O��Z�*h�!Pm��{)���"OnT)�mQ7TJ�=��S�4:|�"Ot���(Y�N�����eZ�R��(�"Op��"�S�_�l����!�Nd�E"O���儂���q@〱}��dZ�"O��r-IK@�o]�	�C��y�E���@� ��]daCL_1�y�GۏN:v$c��F:����N��y�@S{��rщ�sJ�)s�)���y/mi�}���P?h6��ED0�ybɑ�w���HC��#k ��`J���yr�� 1[�h�s��)�N��U/B;�y�I��wS�qR�W�?�p�$��y�f��dln���$�?{u
����[��yR�=3��hP��5w)p�� N��yR��'	��(�cM�y��˩o���"�N�3B���yI=�V�j�E�,)�d�I߯ݰ?�K(#x�!�@E�%rWP��x:��y��:4�� `"�Ė 6y��Y!?�飃�I&Mf�q!�w�'}��0;�
Ҙa��xa�o��xn���=z�H�7�B��Ȱ�L=��zA$l@�n�I��ҧ��d�adaոKn-����`n�t�S"O��2�&H�X<�x�P;AE2�3��p�����s��|�G�' ^$Bv�ڢ[��dB6����T��hb$Uc1��0n�[u$ 4%�N0[�a��#��Y�	0�42҅�$>�p}YG�
Qg�l�b	.�GC�x�4��,,���>	�7FV��f� �n)�2�K &B��!S�H��C߶$70����<���	�(=�]+�Cұ�S�Oפ�(�G�	|1�,S�F�����':���J;%�ʗ�?]:���O�-4�޽t�`��Wd^uի�;Vʘ-���
ن�I�r�x�B3ꚃjh��0q�Ю9@q���ٷ0�4$��
On,�E$7 �@*ίx�D���I�'T���D���"q��9�� w`�p�4�ʨ�����"O��%��1GV*q�QA̚z�r�'0O�[E�Τ�O��%/9.�%� ��)�)Y��@�6q�SJ-D�l�V�4*l��)Cb:Pܹ(}BƄ�w)&��#G^P�ɉv-,��cW?Y�g+�T���'�%>�8��i&�O4Š��ּ15���G�@|�4�	�#�Kl��(3<��	���`�!��x�K�	12���҃*)�	Cvn���x��f�D��fæF�LIHP� �X�:0!6Uni>d��I�V`R$qD�z�<�7� c�\���Ш���L?��D0I%�l2�[�`�\�&�
-j!��Յr��ܲ�KE�8��y�h,`�'s�)�3��;]ʴF�T!MX� `i$�����Β�y�I�,��5k��Kw:"���b�,
L�(࢞>1�IE_���'-BWc�x�	��(��7ܨi��'ȡ�"�B�Ĺ���3~\�RF�;e'��y�Kx�`�DA\(]8������K�AT��ay�cJ:4�(2'i�da\j�~�ؕ����lB�A��4(�B�I��b�{���/c�Ȁ)�n�F2hO
�1�`\(S�h�x�a�u
0����aθ0�j@����6ne�5����?i�!N�1;6���`R�;g��A�@�bټ�����i,=���9V@9�۟	94b>O�ع0� r_t	p���
�f1�a���x�����c�'y�B�@��ڼ �����cG�\����4�ԋV��0���[4b���>,O�A���R�l���f�A�XG��	��O@m�%`ĶP
0�2J����	o�|�U�ɜ%��qвl_{��|�1C[�A�r&#���}�ē%�s@m�tw��2Ŧ"ր��O�l����'A���  t����.}"7��!
u�[���c��+ ��er��'����F��.{����䇾Q���)�B4[W�!�7)N�_Gj�{�LOP*��h�~�(�Y�yR�))�%���A���3�s��M��E!_�b>���-��d�#� )��T��o�<�ӭԌa��p	*,O������~M���pD����O��T��s��3J���TDkݐ����� ?-�p� ҆[��Ri�N>��x�CT>z�b�ᬊ��,�z����w-dq�U.�d~���l��|�O^LQk d��|��\0#�&r��

��j��`	5MA�#4��(�pz�p�D�n�dL�b�1�����,�)ڧDv���&G9~�q2��0#�F~���7<���S���%����@�+iBH��&��!��g�6��ЎޟpF�U{�ā8`�	;{}��G�哒x�����:.����(T(�B�I$	Bp���z�hL�Ɗ��вB�I��=�`�ƫq�f�hGg
>l�vC�87�<�+""�%|�S�J @w:�c��û# �P*O������O2 (�!
!�T@��E\KB�'	�j�肃jH��݊{�@�$'g�ez�Ӑ;�ޥ���1yb��A��Ν��x��E^����jW#;Q��-�~bF�n�ԉs�Ȏ�?Uӳ���z&nDʶ�Ͽ��Y�-�h=�N�?dNd���)v�<��Hىc�V]��HD?��eiE .>���pj$z�L�K�ݔSJ��z%�'�擁V���4��x�D*c6¥b�e�z��{rc+u\���Ǭ�ަ9��jJ1�����ɑ6�|�P7&��.��(�p�
����W�vi*8�Ҋ�3�HO&M(���!Wc��P��4i&��՜%��e���ϊ�?!��S>�F�Q����� 8 *3c�1#�l����q�$ã7?�,c�kAFX����@,W���r�J��*�$	=|��I��?���P�E���G������K��:�di�A��ó+LHqv)"��Ak&D�@�Y7�L��b�YQ�r���2�Ak�E�/���ԫ���aL �g��C1���dB�iھ��{v@�x�t8K�ҔT��P@������=YUn��Б!  z�N��"g�)t�<�m�æq�Ɨ� Nx�s	ԻP�й����M�2�w�;�B7�8���)܆�~��˰�x%��
�$��Wlɮ�y�����T�~���J7�ʲ�|�S� ��,�n���T�:]�����ņ *�D�q'Ƶ;B%���
�M�0��k?�؀V��(�O(H��ϼp�n=�@Дl�ܥ����5[���;�ꖢhYɶ�ݚ�,L�'U�M;P��?��@�0v��Q����=�P���AW��@2g͟��2Շ�I�9�<M��>.��<!pFPG�6��e�	:��X�o�g Y�̓>Y�©�������CO�d�W�%q��l���J; wr���'4�������5G\Y�N��yrȓid�d�S�Ӕ �q��
����q�( |�{`��3���p��[±�r`�}y��l�I���R�Nn��%vk�dm��^���I���.M.�\1ѵ��`���-��K��5����vu���W`L%!	h�c��'S��y/O�0�K�n���qO씢g�U�~����_9N�ђ1�(yqR��'m��oL졛p�.5�Χ����d޻K��9��񉱎�O�n��@�* �#���ܙ��j�^X�"DeG5G7֥/��Œ���I0RR� ѐ�_1A�:QA�Y�J�$e���=s$��HS6�G� �JA�#$�<)M>}ܔ��}%fx
��%C�LXFzBB�	0��Y�oZ��q"�&E�XD*�&�z�4���aع)�~�����Sj򐁧B*,����n�OZ ��/}be=�S9R�ޕX��F=}��D����P8�6�];�ĐǏ�M�R���1�P�C"��E����-F�s��*vk�Ent�l�n��dk'@
/��n��l{ *�3�$Ҵ3�,��"�ߡF���$C(Qk�MÛ*���!L.rX��qBd�t�o�!bx�����y�)�b�P�Cc�D���f̖��0?9F]Lk+㏍;���j�K�J�$�� �5�ؐ#��C���T�i���'sў�:3��Zr qpҤ�t�"M�'|O��iG��Fr�2۴KB}B�-Ԇn�$���GM"T�dT'U�Fi��	�M� x;�� -�(z&�:�l"<I��ڌ�BI���)Q؜��	Z=Cl�}�4r�-��O�*��w�/��䈓�݂<��	�풊z�4��=E��d�P�0 ����eF)D�A#(D�ȥ�PL�d��CGÚad��Y'%3D��2��@�΄�vO�X��qe=D� 9c��T8왅$n�=5A$D���a�
0*���@��)�e�6�$D�`��˨z�xP���-�����y�(E�i|�yp��r�~��
͔�y��%>H�"U�Äj� `bsL�-�yB��Kp�@ƃX�X��͒�y��F�Bd��Iᣄ�'��J��y�d&~���E��n������ybϕ�ZD�v�ޒ	RT5r�@@�y�+�Q��T��_3q���Y�O��y�0k�ԙr�L�e���0��N��yA��x�N��F� QNz��M��y�g�"T���@Y��];f�ȇ� D�tO�9ؐ$r�\��j�X�2D��[��H�l�i3`��V�X�d�.D���'�jj�
�2g����0D�����&"��Y�'g^�D�Ųa`/D�0�4K�	�� �`K��C޲���K>D�$K��B�1ʹsT���h�8t:D����N�J#ƭ�-9Ulu�a6D��k��[�Gc���#X+~����u�6D�<Q��"��!f	HM��;d@2D�D�U��H� �#/�Iq���`2D�\���'-l�Z� 
�"6,��Ӎ/D��3��_;vQ��RW\0
���-D�K2�c�b��	ѾLZA���)D�$Sч����9{�OZ�T9bv�9D��C`��s�HL��� o����#D�P��A�~%t(�׍(��8��� D��Xe&\0hB��P?��l3q ?D���vO�6�f�n��y0�TS�=D�� �+����`��u���U�"OR�!�m�(-� �!�5>�<t)�"O�xHw�]�%�}�c��aK�!�a"Oʹ[�	��0�Ɍ9ԩ�D"O^�B�M/Op>��'�>p<��`�"O�]P�-�h�@�"�hJ�C:��u"O1�G#�0Z]2a�
\80T`�"O�Q��e����5��D~yh0"ObRpGבP� p�. 5,����"O��b���'])6�c���S1hЁ"O�]x�9M��t��Mů)W���"O��14��$V5��A�]�@��!"OD�XHJ4j!h� ��	|�h��"O^�{"k��c2n��K\�'X��"O Y	1J�_n�dj�*ӂ �b"O��S�Dhi�� z$�	�"Oؘ���J-/G��4��4cVER"O����"ܚa8p��'@ԥ4CXE�1"O��ɗ��Pr��2� 5��#1"O<ك���A9rY8�N�a��!�"OJUq��K���1Z��]�w"OhH�gk�8ZK��y�cU��D���"O�蘁ˁ�HH6��:�=@�"O��إn		g��9�K�J.�E��"O��R"��GC� Ò`Y�K���X�"O��	w��Z	Z���%
���U�'�����;tv`P�nD�WfZDœ�L��|��'m��%	X>yɄ��0D��'.�� VgC�8}+���"����'�VH��B�_��	�Z��'{ ��&�ĞAWty�U�F�(ި���'��Mr�!�<!�~�kei��$�,�Z�'~��!%� ,z�S�O���
�'�d*���,("t8e썉#��	;�'�<}� #�(4~8k�bΈ��$x�'�ݒ����6<n����o���'�eK`�Ő{�@a�En�=.���'"N�����;p�x��-�6�2���'X:U��D� �rD5�+��D��'�x�C���=F���$�,�(\J�'������$J�s��ܓ�8��'3��Y���Z���{EI��
=�	�'ovq"Ѓ�
@:�� J��/� P�yb�5�ŞK�� �)�#C�`�d�Ǐ'Ap��'��A��ԟ&I�I�PB�JWm��!�p̚�%-6���p�T���MS1���h���ݘ2 A����	
BDP�F�#2p�i`�e�0t�S}�O6�u;F��W�T��+[�&�b�q#�$S�`���~���y"g�f>}�T��:7�����Z�y�A3~2	S���*��,"1J�'�y�Lϖj_���&��\�`�ݎ�y���:$��Ή��у �2�y�T<P p  ��   �  S  �  i  h)  x4  f?  �J  %V  �a  �k  &t  {  I�  G�  ��  �  8�  z�  ��  ��  Z�  ��  �  k�  ��  9�  ��  �  Y�  ��  c�    a � � � ' �/ �5  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z�����W��K�L12$���SO�\1Yd�	�O�!�WR�H�Ī�.b�&hb1[��Q�|���T>�%		i�JI����z�`��6#1D��Sea�d]`b%�\th35D������?!�-Q�ė
?<��F.D�@3A�	5�Fy�B@WD&�H�!D�,s���CB>�rR�>dwA�*D�$0R�Ō*���B��30�)�-&D� c3�jFM �jp����('�ب�^��*�\�Xi��tU<Z "OlA�g`�$`&�@��I�kHH\C#�'ў�
Q�� P���]>�h���$D�\��.�h���p h�X�\�L-D������~`&A��K 1.V���5D�x�`ך_s��:��Yd8�4?ю��S7\�^5 A�ݯ�R=8�'��B�IP�&D���� �DU� �#$��B�I*1	@��G���J$E��LOO�JC�ɨp�\Dhfe�?`��鱺@�e��=O��i��b�x�Y�)[�ks$�ȓk��b#͔)rNQ��K�j>-����@�w�B�[*�� G<@�-�����DNA�R}�U�$���g\�܇��i��T}���.Ƞ��ĩ�C�(��C�	\?ы��?vԠ�F��K�#=���T?t���N�\Ry��:D��ۢ�b0t1��,�'b�tg8D����d�M{��CK,h�����5D�g�7Zr�#�o�!}�%3�B4D�pn\t���V͞؎i�sG0D��ڀK��/��r"�0�r%)��.D���u#�l<���`��MfNݲ�M-D�J���p���s�mX�1F�K7,D�PsC�Rj�����RLmXB%D�d�5mc�D��aiT�u:8}��#D�Da�H/6)bY�dݹV(Yxu�-D��Ԇۜ��e+���
Z�H�c+D��c[1N��A���5���R�j-D�xJ��S�u����@�b�``���,��h�4`Gf����B�f��C�Y�h �ȓ&4e�R�:�t�Bt���4!�ȓiW��
G��#�>L�s��)�z��ȓ3��Ց�B�	N)��ܞ.�4���o\\x��63X�p!Q��2����r��)9V	�4!(�E��
yI0��ȓN#�S ���(HG�ϭs�b�ȓM�@�y��/^��6"L�Q�ȓT��"��԰�h���֡�X��gX����H��O \�j��%g��ȓ.��0r��ݍ4�8�Q�<o]
@��I�L�Ӄ	"&^B���ǻ)�r���<�@,h"�L�\.t�%��6���+݆=s3��W���!DK҅��݄ȓ�z(��k���V��EU�j0���ȓ�R�Z��L�^��+��Q�k2(�g��~b��Y2���Mۉ\�����[��Ov�'	|�c)�*P�ӋA�1��Tr��,|]
g"O� t��v��,l��A�i�#�A�R_����)ҧ �`gc��Qq��a�.Jž�ȓT��1ٶKW Ĥ��@Ж3[^�%��z �'���W��-�:P�gK�.�p�'��Vhe����ȝ����9�bB�ɚC'B$XEi�3Q���R�( ����RO�tJ��BЅV�h�k�$G�n���BG(�<J��C;c��Ӳb[7L��09s*LO7/�I�QT�b�-��,r^ѳ'ɍ3?�*B�ɕ{�z�12LD�|��x9r�e�RC�I�f7�a��`� }�D�����B�I�5cZ����P9��S"S�84�"<�:��A�����Hy>���M�9#.�@�ȓC|��+t�/)<e@C��7hL�ȓ~��)��X9{���R��;'�<ф�J��,E�F)�prc��r���ȓ&e��[���88�£�8Mu�q�ȓ]o���1(�v�z���0rp���S��,�?W�Rqj��0)���ȓv�
�p��<@��x�t�������{Q����nU{��@�FF�����J���7 J%M��1)P ԂC�Fź]�� �5ݺ vNQ�a]�C�	(,�x�H �+��PC0!�)O�xC�I�$ޔreM�]J�s�OO�%�C�I��
��
�;.b��Q�����@B�	�Sh�H U��2d��vޟwu�C�ɐE������ ,B�2aA��j2xC䉏*hTŁw���x�ʴ�Z�}NC�	=<a��j�#9ZB [,W*�<C�I/odٚ&KиO��32j�>C��妰pb�S<(�6���'���e��&Pb���+ƾi�0ES���|m���Di6ʄD44$�[�oI0�^���>͌�*R���+�,�$%`��&v��Y�G�D���\�kڦĆȓ?8��(p�-^`<E�.��d��,��2B�ܻA������=��ȓq�*M30a B��r�
Ѭ��ȓ4ᐥ�$�G� ��u�s�x�\͇� xp� !�\��Ӆ�f����\6����?O����L��$�\�����I?e����$BXQc"O0�t��~�����L1}0��{�"Of�����x_y�3mυn(D���"O��ue� .��AQĂGT�c�"O�к%'��_�� (��N�;�>-)�"OT%���N=$��0f1=�Zغf"O�3�ɒ�}��%E��_��5"O ��g̓��V}X��ܖu|�1�v"O��h3�Ɨ$b(+����'U�)�"O���p��E�P0���s6�hA "O���1���!?@P��ͽ[���"OH�	c�$z���q��W�hXX� �"O�,�!FL��`@� ˭0@��"O���H��"�:�po��>:�""O&�h���Uc@��w/�uS�"O�9���N0�@V�r p�0�"O�K�b�g���9WE����	�"O��@��˜txs��u���:�"O*���e�j&ਣq�Ʌ:�xa�"O�X#`gE� & H�%�S���:�'�u�aL�ބ	������6D��2�gX�Fl�!�fG�5N��e)3D�� xk��+�:��Ç�'���d"Of%k�߃3s�l��On���"O�0;r��(A0E#�Í�5VΜ��"O��炍S��(� ��Er��J�"O�첗������*ݜA�Z-���'3��'���'b�'2�'�"�'=Ҹ���O�:�
9��pxF51��'V��'���'I2�'���'B�'X�)�w˗�c��] �Λ�c5��0B�'���'��'	��'���'}B�'���[���,8xT�,ݎjڌ�4�'R�'�B�'qb�'.r�':��'}��[ 
жO>^ԋ�6	��P#�'�2�'�B�'5R�'��'���'�0T��ˎ�uW��a�h]�0�4=���'���'���'b�',��'�"�'��\���l��Fj��JM��':2�'��'��'��'���'�]C@��'k�����^;P�����'9�'���'T��'H�'���'QlpZ�D���'���l1��'"�'�r�'+��'��'�b�'x�U�As}�IE���Z����'j�'ob�'��'k"�'�2�'d�ū� K;6\d�C�[�aNİ�e�'4��'���'!�' "�'D��':43׮�Q���jҋ�"dR����'�2�'�r�'jr�'���'Xr�'�8�[W�+&WV}c��C�H0��'���'-�'{��'���b�J���O4�I�;'� )��ܒW�L	geCy�'J�)�3?��i��M#Q$߼P�\�8T��4p+��۝'D�	�M�R��>��@$�m(E
,�$���Ŵa ���?�,Η�M��O�瓸�rI?��v��'O�L8��ޚdJ�v)�ڟ�'��>�3��	 ~��,�&�8.%�r��4��D�<����O0�6=�fQ���&mD�S%ʟ9�|�1fh�O��D|�pԧ�O��}@Ĳi��d��o����G[��H��D�<U��|��� �L�=�'�?��S�:��7䞘MA 
VHL�<)O4�O"��~z��C�8����Pol��d��m�<i�2N�>����?�'�I�h����!k�%��ѹ��ΦBx��?Aԡ
D�:l�|Bā�O8l"�n������G҉��Q���:(O˓�?E��'�Q15�QC-n0�f���*���'hd���D���?�;Hm�5��$&ZLɊ�o׷z���Γ�?a��:m�%
�n�j~�:�����F�4|I������G�ҙY��!&�|[�b>c�(���Xi,�򵆞>�2	�f+?�X��� �Ij��/ڹ��<�F�Kg�K�aL1SQ���Iڟ�$�b>�����v��*HQ�u�VNSϒ�`�ISy�i�/9H!��%UE�'8�I�{B�0�S�\�LQ��@Ż[�T�����	��i>��'����?��T�B�~Yʦ�  &px�BN��?��i��O=�'���'2�R�l𙔇݂t7H�c'9G� 6�i��	�!��0˵���U���+�ҵXC�?��XwBr������r܀����]'ۂ,{#�R���h�	���I����?��4��L(3�K-\S�1�٨H>��?�'QyA{�4����(S�	y��4��Iɋ���v��~ݞ��O�����D�OL���O���E"�p�␋G�-�f�20��\e��d�O�����������x�O�u���ʧ{U��e`
�a�h1��O�@�'���'jɧ�I�l3Hi��� �ֹ�"fS!c3Ơ�4#w��v�2�����jl?QO>h
�u�lE��CΤ�����F��?!��?	���?�|Z+O&�nZ���d��=Z�*��&.�\�.�	`y�mx��⟄��O*���'*f�I#Cɞ�r��	Ȫc�����O�;&t�t�ҠP�w��>�O<�T�sd˾@�$�5�ƄQ��d�'C��$��ڟ��I�H��k��fI�d4��*�%���0m_���?����?yK~��JV��w�����gӆ�a�B&4���"�'���|��H %�6>Ot�)�ݼd��͡��]�GoP�R:O�����?)�&5�Ľ<ͧ�?y&�^�2��Aϳ9^9������?���?!���dXp}r�'���':DݫSO��q����u'��	b%"��h}R�'��|�k�=-��b��GT��+�������9���K��wӞc>Q���Ov�D��:�:�#\?�
�#PÔ�p����O���O��?�'�?i�)׿l$P�(�>���+Sѣ�?YR���I؟Pk�4���y��V�\u���6I���1{�T9�yR�'���'0�d;q�i��ɪ}��<ޟ�l�  _�_�@���-="�j�F(�$�<���?A��?	��?��V�����b�$�M�ug<���B}�[����U�̟DˀI��r֦	���ū<T� ���:��D�O��9��I�_�8�ba$^�9_
�TBG3Y�Q"-@+a�Ɏf6��p�',��'��'�Ҍ�2lK�h�q��dϤtܼU��'�Z:���'��O��I����O�|b���+� ���i�^-����O&l�A�U�	˟��i޹��EFBF��SPqR�JrCRz��lla~b+�I��d����'ֿ� �%I��?���H"��8zBݙ�=O����O���O ��O �?ّ⨐�k��KQ���y����ܟ8�	��i�O�S4�M[J>	Q�̨<���h�ǘ"	���ȟ�䓒?��|:���M#�O@T!1j�3'\i�R	��wH)3��nd�9S�'1�'��	̟T��ܟp��M�L(�ç,,Kv�E@Ц,��9�IԟЗ'����?����?�,��٩���|��A�҄���)�'�<)���I��p��q�)*�jC5]��3U� '��9�k�"��TcF�-�M;eT�擶2T��)��rvq.���R<��(�}e�]����?)��?�S�'��T˦i�7eZ�L�J��s��"60|�9��`���I���۴��'����?��֕%ne�d���c�d�6�ͤ�?���#\���4��DG�{Y��O��	 ��ݱ4�N�;(:l��"�7uC��\y��'���'f��'�b^>�(R.�?u/���
���D ˂����O2���Ov��4�DX�����X�%ϧ?�J���E
B�8a���t&�b>��"Oצ��J7X���1ր��FAP�`�ʸ͓\|�A�C��O5@N>�+O����O�$H�6>m�qvN����<j���O����O2�d�<�F^�p��ȟ�	+1�pX ��%��7KÜ��?)wX�p�	�,&������q�ʃ�O�|��1�0�8?9�S�_���z�4q��O����?�`���2��t.�0:�*�c��?����?���?a����O�t�e�
2�;Ъ�8U��)	�#�O�8�'6�	�Mˊ�w\�m��o�o��h�e	��H�'��'Y�CZ0Mܛ���`� ��4&��ۂm ZM�0D�������J�$�)$�������'��'|"�'���r'�q	>��7�'�$}��Y���O����O��!�9O,��F��윁P@5����j�F}b�'��|����?>�MÀ��.� ��.�Dj@�Իi?�	� 0�1�OҒOʓ@TL����3���%ۥ9� <��?���?��|+O��'32��%X8�⡩�$_�bh�O֓¦a�8�T�O�$�O �$A�6��\���MP���`�I�T50]s +l�V�'�����K�n0�O~j�;^�=k@��4u������]����?���?	���?�����O�,�V,P��E�p��������'b�':��|:��q�f�|2AT�Y&lBA^���$��mU8&�'�����T=3�f��H� F�#��U*�CQ�N���A��6�3��'4�&������'0b�'P�M!WNU$�R��VhZ� =F���'��_�0�O����O���|2�)�/�%B4C�>���mY~K�>���?�J>�O�t�rJS*D�����u����JW '1
��"�i��i>� P�O��Ov]`�,����`qLչB�� ��O����O��$�O1�|�E)�o�	�VM�f�� `�ʭ�%- �y�^�P��4��'����?�`D�>�. #di� 9�L�U���?��_=B���4������]��ڙj�!��$�v�!p��T��y�X�������� �Iϟ8�O�D�Q�/%}>�3��N3U��{E�>���?�����?ac��y�*��xu�_�{���W
�F�2���.}�7Mu�$�AD���tYq��7i��;�cj���펔r��|��Uy"�'�beP"J-p�1��w�,H��@L)i��'�b�'5�I��D�Od���O�kt�ϾDĵun�-oBxt�c�-�I����O��$4���=\Y���Aѱ4w�sĄ�2'��	�c3�k@��eD�U'?�{0�'N�q�I+�T ���;[m�8�QHޞ������L�	����G�OC
':BE�L"w����/�Ba�>����?)W�i�O�NÜi�u; dR�O�6�y�-G :��d�Of�$�O��HR�fӜ�Ӻ���Š�J�&A�NH��WG�2���"�L  �O�˓�?����?����?��˘����n��$heM��R�DZ*O�=�'���'}B��ɍ;g�l��6��,�J�(w���'���'Pɧ�O�\5+0cB$�$4�QF�=1��	�FJ�z�º<��lD(<S���w��^y2�ƁD٥.��kP�`Yb�'�b�'��O�ɍ����Oޘ�sH߅ZFA��nG0\c��a��O�l�i��x�����'��(11�����a���&0KZ�X'�ɤ1����(i5`��;O�$�Er���)´A�	W05`7B�.0���c��y���ğ0�	�����֟���@�q.�H�7�}_�"�2�?	���?IV����ٴ������ˑ-��p���P���I>���?�'`XX�۴���?_����h�.|�	�b@�kcXQÖiC��~��|�Q���Iğt�	ß�*b7� h��-CzLŐt
�<��Zy��>a.Oh�D�|��LA�&.��!!=NL�q�W~b`�>���?)J>�OȌ٘��Řn�Y����Xܶ4�̘���-J�'��4��%{�KTv�O��vj��	��C�. 6���f��O����O���O1�j˓|���kA!q'R\
�jv�Xi�ФP��y2�'��wӖ⟜c�Or�Ė�&��ĉB⑏!�N�A���_Gl���Oze���r��Ӻ[@b��¤<� N�I�E��=�2ħ�2?/�I%4O^��?����?����?�����)LK~N�(�M'$]�$���1����'h�'b����'>�6=�\���/P�,�rOA��D+���O���(��i��r�6�i� ��Vg
|tزE��$3�� ��k�q�G�,\�C�J�IBy��'��өO fY�j>� v�TrVR�'�B�'��	����O��D�O�����M� �*�+ ��]ڦ�!�I=���O��$=�D�3]���(R�=��-��Kd��I�7N�Yz�AT$�Nc>ur��'�N��I&G�|k�E�=L��-݄j`��⟠�	̟ �Is�O�bf[�e �����!O*�(HN!ej!�>I��?���i�O��hZi�p�Òhcj�3�jXd���O<���O�<�P�nӞ��$�b�����q�<ߨ]��V�Y��&W�����4����OT���O@�D�,��̑R�ã!�k���_X�ʓ���ٟd�	ןt$?a�	�BŉW�i3!�)yW��٨O����O��O1�� hukU~X	�*��F`�嫂+"�|�����J#��WA�*�A�I@y"J_��I����{���5�n���'��'��O��ɛ����O�a�ą���i��T*Ŭ�y��O4�ow�������������1�W%����i�;3�,�B�o��m�\~���Q�t�Ӌ*#�O����m0�M�0k�[�Kò�y�'�r�'��'*���T	�RECU�O����S!i@���O���`}�O�Bf�֒Of)��,�j`J��
�).T�F��Oʓ5��ܴ��D��0�ڜbC*��=�w
�*��(L��?��@=��<Y��?����?i�?u���9E�X%S��m�e�Q��?�����~}��'���'��/Ia�ݙ�-F��;T풦���2���Οp��\�)׏P�&�di �@�#_�x�y��Ȩp��5��"l����dٟ(I��E�9��(��DB�ݡ3��1CWb�'�2�'<���Z����4^ ���O�(#�M���p�)ϓ�?��M���$W}��'*��"��R*.��m����J�j����'I�?r�6����<.��q�SJ���"�F��Ƨ�+!7���+#��IJy��'���'|��'��_>Ep�ᚖ��D�����Ϯd��)��D�OH�D�O4����ڦ���(��ĵ#�dA*�M3#�r���ӟ|'�b>�;�����y̓=q�����6	��Z�Kr��T̓|��;�`���'�����$�'8��ԯ����AYa�M�i����'���'�RU�TۨO����O��DW�Yi�)�"�="b$�D�dz�Ot��D}��'��|*��0}sp�_�,>�:������T�	j��c҉8IR��J����=I@�$W-�iAI�V��|٣B�w*X���O���O���>ڧ�?y%�R^8�К�ϹvH^}�GϺ�?	dP���'��6�1�i��0S�Z%1�:��&H�U@�T(z����ҟ ��-I��lZ|~�d����k�RM���;`�p����@��|�^��̟��	��	���1!���l�B V2�FXkՍKUy�ʬ>���?�����<��B�&����R�K�� �F��u8��Ɵ\��v�)� -ґW��ZK�Ӛ5_���M��	�'j��94.�D?�J>9/O.-�A#��y-����߰jj!����O�D�O���O�i�<��_�P�iUa3�C�B,6�YSD� )��R�'V6m%������O��$�O� (l\�W\�hs+9W�@� �K�:7m/?	�J8;���4���}�#��8B8c5'F4��1D�l�I����ȟ��	����:�fȁb�\���,�#85��B�������O�,ԧ�d�'j�7-(���4C��p�ǀǈ2�z�:U(��'�P��Pn�����'�����JX�z��̠W�
T�D)��eʠ ����z�'��Iǟ����ɞn��d�G�ӽ5V0���ƈ�
d���	����'oV���d�O��'K��`�&�BE'ܭ
CA_Y��'�l��?�����S�d_�k�� �&@�T9QdF?9t�]�&CڶDLR@:�_���h����|�	�+�u���%�-�"�%/T����Ɵ4�	��H�)��dy!g�j����eo�p�%
,O�N���5Ox�d�On�nH�	ܟt��O�����B\��k�"˄0��T���vL���O��8�`���Ӻ���I����<�ƊX+z�:Y��@�,b6Nd�Sm��<�/O��$�O
��O����ORʧw�ڰ��K3]l,���+F�p�Y���Işl��x�ş�����S�Κ�^�p6�1vN�����:�?9���Ş/���4�yBW�Vgzq[�@���K�d�R�'ez`p���՟KƘ|�T�4�	ß�[��w���0TaS����*լ������ß���ay� �>�-O��d�u��\����m�* ��L��l�t��O���O.�O��`DM�f���AT�E3J|�����ċ#�L�O�\��W�S�H�՟�1� D�p[t㉤Qh�u2�KD؟��	�p�I���D���'�x��%�#���a�������'mN듺?���r���4�*� �h 2Wb�k�"�h ���?OF�$�O��䙋h�65?A«�l�����c�? D0�E�Sb�L�"e�?0 �Ղ�c$�d�<ͧ�?9���?)��?�Q˚
��̢`�M$�zYH��А��v}��'|��'�O~�-�"k�F�Ч(�����K��p��?A�����Ir"@�d.��%rQ��@w�qq#B�Y��	L �q��'Pf]'���'�,��&�Rfv�ɗ�1j�]ʣ�'�'A���dT��	�Ob��ƙKv�I��3}��	J2�]	Nbj�$ܦ��?�V������ɪ,M؀*%�1(~�q㖠=ob� �MDɦ��'����E
�S�O�w��t:Թ�D:|�vr��B��yr�'Qb�'�2�'��)Lo��A�m>��d�eg������O����y}�O��%}Ӓ�O\YC�E�g5���c��{�nf�5�d�O��4�)3�d�,�Ӻ��%ڐI�xk��o�L<*v��,�����c1̒O�˓�?9���?!�J9��C��ri��@H�⩢��?�(OBq�'RR�'w"Y>�ٱΰ��%A"�I/Vd=�k3?��U�<�	��'��'0����^-G���y�H��1������'4a3v��R~�OZ*|��%��'y�E�a�C�lv���y�8k��'."�'F2���O�	�M�@i]�E� �o4� ��L�<A���?Q�i��O6��'T��Q5Xܸ;%��<d�°�s�S)�'��X�d�i^�I7�N�b�	U�x/,尶b�C���st��"l5�<����?���?a���?(����$]�}�|�{]��嗦$
�P�':��'�B����'�7=�\p "�9�훇�үt?�����O"�b>ͰB˦͓UuP��`m�G�L��4��O�j�̓
֚��i�O,�L>),O,�$�O@ ss�޹:gJQ*Wa�555~Y�"�O����O��<��]�,���t�I�}$����,kСK�d�GD��?y�S���	ܟ�'��+Ǖ ��)�o]v���%$?A4Dպ+�,e
�A�'#�&�D��?�U���b��1CV��8.�d��d�U��?���?����?���i�O�D���K%~� �጑�F���c�OЬ�'��'\ 6�-�D�O�F0X�*(a�N�Ig�i3En�.v���On���OjѰ +i�,�Ӻ�G�Y���K�~V��aL�U� �V*kv�O���?����?���?!�a{�c��I.?�a����13�Y�,O*�'eR�'GR��t�'��<s�aXY�
)�i�l	��!�>����?	H>�|�b��L ����Y�x��8��	/�
���4���W�0�~(3�'��';�	�+$���z�:A(�M�a������Iϟ��i>q�'6듥?�%	V`IF�wO���4�����0�?���i��O�%�'���'��G�gSؘ�� 2�`���ɺOd$%�id�I$�>�Y�Olq���Nҡ:B��9v�G�0?��
!�R(��D�O ���Ot�$�O���-��"0X��La�H\�2.�?Q���ß����4�������$��#�0�:��ês,^١3��|������i>%��W����'�d�C��\(�J�h�+q�$���,^uʕ�I�F�'v�i>�I̟����.!p	���[�2�x41�G��x�t=��ПD�'Ϟ�����O��'^A&�(UF�6g�a"	�6�ı�'����?�ʟ���gߚ\�.�@�,e�d�A�OgFV$�p�&���|��Ob�O>A5�A5n��XYҧ�&��|����?Q��?����?�|:+O25n�2�����ƶJ�hY���B"��IXy�Fw��DY�Op�d��V=��bhS�{A�qa c�П����*eo�z~"ꑱ��}�1,��5�p8D�$@
h��#�<q+O~�$�O����O����OZ�'UnXpEU.�v�R�7Wd幰V�`�'b��$�'V�6��l�:Р���L" ��#��'	"�|���o�8r�64O�1H���.fP��!��;%�<��;O.����?�S�,�D�<1+Ojh���!-O(\!�Բq� +a�'�r��?���?���@W�	���Q��p�o�'��'��듐?�������,���|�8,s�kL+3�DT�'��Yf��D2��w��d��ݟ����']f%E�PTj@aEj�.C���'�b�'�R�'a�>}�I�HDT��R��`�nM��ʓ�q ��I7���O���
�}�?�;�B�PulކkP����+s[@M��?����?)e�K'�M[�O0i��*��Z�"J�(�v�ۑ��Y�Bxz� ��m��OD��|����?I��?��i�ȹ��	ƀ��@�P)F�(F^m�,O8|�'U�	ܟ�$?Q����Q��L�-S�A5��s�O��>�)��6������_*ʉ@��D��Ѥ�Į(�䨕'�����ßD�3�|�W���#*�,N��D��lY����U�۟��	��I��}y�>a��|�h�%�	�k��,�u-��Q=��+��Es�&�D�X}��'#�	5L<�@ӒI3�&� ���D��Dґ��ᦽ�'W�
�MS�?q@R��$�w���J�#�%s|�X0���k�8Ź�'>"�'lr�'��'/�P}��A�$@@���I�L� 9tB�<a��?��i>9�I��M�K>b��%g��`"3-�P �q�!���?���|b��S��M��O�+p� Dh2��	q�.5��%ʳ,�F%��Ʀ�?A��2�Ħ<�'�?����?�ס�>}�����>10�B�J�?i����^}��' r�']��K[�< ��9H�:l�B�����n����� �?�O�>@)V��0��bBD�W���냙bbT�q���8.�i>�A�'�$�<�$lم&�h
T�A&�<ᒆ������쟔�	�b>�'�Z7�V=+ �تU�Y$\k�4zB�S��$�O���
�Y�?a�X�\�ɣX�"Ę�΅-rOrMr@㎵$���I͟�!5-��A�'7f�r!���?������#�Z�Bcz,k�o	�j��t1O���?9���?����?A�����	�7����áLh���E�H�'�'�b���'��6=�b�ڥ���l0��+��ݙ%�x��/�Ox��/��	јɬ6�{� � ��!�y��7blxpz��Y�v�"!�D�I[y2�'OR��6@�j����;yx@4�M��2B�'nr�'��I�����O���O2��p��\&NY��ļ
�^���2�������ON��%�D�|z�報ʛ;5��ʐO�|���7w^�Uq��\9�c>ay��'�M�Id�.��wɉ�#� E	��9F����Ο��������G�OM�FE�R�z5C��8b�Qf��$g�n�>���?���i��O�P�\ iBf�8kz�H��Y91���O���OV�K�,{�j�2���Fά?�)Ǎ��
[�͋*�

�Na�U�Z�	Jy��'���'gR�'$⎐"�����,
$^a�dH5O����ɿ����OF�$�O�����2t���RA{�I�I�Z�:��'�B�'ɧ�O騈R�&(�)���F^�p�7�͍#��v�<���˽8nf�IJ��]yBAE�?�~ԣ�ώ*tp��`,L%"�'�R�'��O��	����O���Do[�v(d�RWM_?i�\p�v��O�QoZM��k���Ο�������$�U.S��C���9/��]��"���4����=�Ra:����O�g�_�~pő���VJ��U�y�'�r�'0��'(2�	���,�.�+��
G��<5k����O���Wf}�Og�$i�z�O�X�r@ιV[�X��O���R�D*���O
�4���1V�t�v�-��p�ˢ[h�4�"PJ�̙r��
!���K��䓠�4�`���O����Rez�۶gX��]�a Ƶ���O2�$�<�^�t�����L�$P��mY�*A-<�ʘ@���y2�'���?���O�"��s���c����0`���zY��Z��	���BpW�`�S�&��_�&z^�i`�'L�V�<���Qxi���Iɟ��	ğ��)��Ky�Jy�hY[��ʆ	�l���C�!UΑ��<O����OT�l�x��	1�	ݟT���J5��:"�͇8�h|�`�Vş\�����m�D~Zw��*R�O�h\�'\P�Q��_�K~�͸"!�����'���ğ�I۟(��ӟ�Ih��K}[z���O��$��`�G�;����?���?qL~Γv	��wN4�iƅ����C��A�~;f;��'2�|���#]�NU�4Ofd���"
����NP�6=�4O�y��A��?Q�O3�D�<ͧ�?1�M�:�x���h!�A�7����?����?����D A}�'���'>f(*!-��iݲ�����	}T@s����N}"�'}��|BcX,���#�O3�L�zGnE��$�*N�����Њ�1�������j��O�6�^ �ІРDe�=����b�X���O����OD��%ڧ�?��䕪'P��Lî|�:��4L��?��Q�����$��4���y��� �q�1V@Z��4jD'�yR�'C��'�}���i&�Ɇ�,���O����O��W�mK��X���L��%}��Oy�O"�'��'��˩X�d�!V�2�� k��J��	��D�O�D�O~����J?�Q��l^> �v%ȳ� \�� �'S��'*ɧ�Oݢ��A�B%7Xn���أT[��kF�Tq,|J�O�����β�?��$+���<��bL9]�օ� ǽ4&�5�!g[�?)��?	���?�'��F}��'����`Ј_�*���i��~6d}C�'$"7�5�I���O,�m�('D��md��dEQ�2y�i����M��O��W��� c:������(iE�@�GJ}�f<+a4O����O����O��$�O��?IB�$�T��vN$A]����䟼�	����O���O�Moh�J�����f� �1�ܔV:8$� ����Sg�2}m�Y~����;�jY`��Г.�j�r�Q��$E�Ќ�ğ�r�|�\������������8E��B�̋v[L�X ����	yy��>���?!���	0K�B�j�jQ�'��c"�"��,��$�O��$%��?�3��W�o�Ds��6j)�1hVc_:#Л�Ɋ��M��O�Ɉ8N�QC��(.���"���I�h1�T"�lT���o�LP�A+D�Ne(F��j�X���k�$��DnV�TxA��+X�Wf퉴�J�o��5`�Yf��aW��-�dٱc��OH�Y2�y�X¥䆍bG�M �e�3m��ce�;�|�1��X���cM4LF0ѢK�Itp -9x�a(B�=?Wp�pf̀;Lhd�Ga�V�+���w��E���,n��ݻ@�R�,���І�Y��@�B�h޺@% �B�B�x=	�Z4_�E����-�-¶昄NrTX���g�4�1�i����$�Of�O���Ox�����Kr���po[Y��x�p��� �dפt���O^��O����3� � q�Q7F�x�)�F� 7��b�i!��'��|��'��,�3 QZc�98!'[�(�s�/ �L���n`���Iʟ �Ɇ��'H`��ǟ<8aO�76KL�KQ�(��\���H��M������?���4s�{B�BZRt��� �m�$�,�Mk��?Q@b]�<a�����O����O��be�BWiZ4�B%Q	/��Ԫ�j�f�	⟬�I)� ]�?�O�f� 2/�~L��F�Jv��k�4l�x̓�?����?����?���$�.V툍�4��L*H�@$$Dq�mZ�p��g<���?�O{M�شp,<I�U��'$�8�@D�␩m��|�ܴ�?1���?q��k���Hy�JR�����?I�K9�p��i8m���d�|�PB�<��U��R֯ޣ�H�����7OgFa!��i���'���'l�����O��I�]� 8�d�H&	7��@�*Q*.�c�,��OG˟���m���۟�	3 F�%�%�U�pn�xR�/z�q��4�?)�vL�IVyB�'�ɧ5֦
^n�9�ïrJ	��I���� �tyr���;2���O����O�O�<�w�̐*W�!9]�Qoߟ�M[�_�4�'���|��'�2f�\zb�O4L�2���Ԑ,��A�'��8�'yB�'Oҕ�dz>��Q/��Eb@�a��0g6�8�k��˓�?�I>��?��Ɂ"�~��t�����E�I&�a������u5O���O��d�P�SX�t�'�ҭ� �`(�� �͔�S�X\1VDe��!���O �� �w��ؓ�n-Zv��EN�e��bhnӂ�d�OT=�B3O �d t���'��5��ɢcRpP��\	�����F	������ON��/�9O�N' 9�Dkc���+���iU"]���˘%�yR�'�7��O~���O*��\p~�ߨm� ��mr�\�5,x	o�hy��'�b�1�i�|.���I�n �B� �3g�PDs�ǆ
%�Iܟ��	՟�Iן�������1�L�f��,��fi�4YN�E�'p��#��4��y���ܙ�a�v�pч3g�*F��6�M��?��?�.O�Sa���'f�S�"V/"ux�kJ�.@Dx"�}�����"?���?��@T�������8� ��__|o�蟐��XyB"�~*��j�)B�^�S��ٲ]�"�k��ǘ5�O�s kR0N������i>	��tغ��#�	
#z�����v��nWyr�'Y2��O�I?A�vM�%��*qJʍ�s�C�,t7�vJ�ɣґ�d�I՟��RyBџ�	�R#ֱ@�*4�æ�"\��ԷiC"�'?�O�ħ<)#hFϦ���)_��prf�*Cxͣ��0�y�'|�'S����OR�)_�*܁J�H?�� 
V�G(��6M�Oz�O@��|�����ʔ1�C� �õ�k7��O����8�\�,�O��'+Zc!�d�cN�tڕ��HƣD�x�K<!����\����]+�� �E�Q�g�J@�d�hp�7mȦA�$�O^�mȟ���$�ɑ��$�o<V,k��v������4T��]����ן�J|r/�.��p�i�6�i��K�@!jp��&&���O���O���O~�ī<�O~4�^aP(@5��?!?T� o�>y��W����!��y�'�q ) �c�Òj�*1ɑ�qӲ���O(���O�<&��'�~r�Y�� hh�)ԁo��L����M������?���<1��2۴�?��KP���G� �$���#؋	���'��n8�?��'�iY�m�dq��� ��Ӥ��5$��',��y��'���'����� ©� ���Kv�F�n��-nچ���?I��䓚��$�!��8�) n�BfP�!p�i
B���yr�'��'*�O�H�ӵ��0�#F�xT�%����ISv��?����䓰�4���d�~��t��@P�aZwM���� 1Op��O�v�Ӊ��i�O�t�!n�>Pr�Ui1ǜ��`�s�B�ɦ���vy�'�2�'��4��O��^�\y:6͂�j��A�T�m�<6m�O��*|��D�O&��O R�'���+#��L��.��.�)���?x����?���?�ǡN�<y���?i�nM�(L���Ϧ=I�Q�|�<Pr�:O��������ş4�	�8!�O�NΗa�mjeNAb��풁j3�&�'�b����y"�|X>�`�tӖ,9S�xX^\p��|�L1�ߤ%^�`k�v��O����O�a�'��ɗ0ȼ8�� !
�2�.��XǨ��޴o��Γ�?�+OX�'=9.��'�?Qp�E.(N�!7d�O]��@�j�DÛv�'���'H�>!/OR�d��$��=��1
���m6L����v�T��<A���<�voP�|
���?��b��PKJ���Ju���~#,PW�iB�'Q�����O�ʓ�?�1;%@��dV������d JM���'ڼY��'����u�'���'����yZwf8���Ӟk~�M`f��
�R�2�4m=��Fy"�'��Ɵ�����;��̏7����q�2b��Z@��7]����'d� �	���Iȟ�%?�ȝO�t�e�3O�ڌ���B'n��)�4��D�O˓�?q���?��'Ha}����E�x��4���h^Ċ�iԴk���I�P�	럴@Yw������Ok��q���R<f��,�%/�F�'��I�|�Iџ�S��(�s�򐚳BW�dJ()��L֩7Ʈ��idR�'bn4��'K�	�~R��?Y��1+� �R֩��Rd�B��]d��2�_�,������	�S�@y��'����na����� �:�$��2˛6��y��'�6��OV�D�O0�\R}ZwL����߹!X�� ���(�:ͨݴ�?1��8=̓�䓒򉙒Y���/�#N����dO�dK6iд��!�M��BZ���'b�'��'�>�(Olq
�
�V;��Qc�W����
��Ҧŀ�h���I^y�P>	��m>���	.N�1 ���c QA$�_ e�2��4�?����?	�3��Wy�'/���Y�0#���3]��͚D�" ��ayb.W�y����4�'�r�'�~Q�K]�{�V&O�]�*IS�(�b�d�O:��'��ޟ8�'�Zc�d�"���	3n]b��Đv|`m�OD���<OxI�D�O>���O@�D���f�����iM��{�� 6G�0h��i/�ꓓ��Ox��?y���?I��R�.��$"�Ex�X�En�(���5݌�ϓ�?!���?�L~�5ܟ<9��Y�?�Va�垦d]T�L<������?����c��#,J��!�p��+�T�8�#��<1���?���\ÉO}|��2�4T��ٯw�|ڣ�����@��i �|��'!��S�yҐ>q�M�k*�򠃔G��M�Un�Ŧ5�Iԟ�k'`��	 ��I�O����O�Tʄ��9�ZyB��I�8.�#TŒC��ӟX��){�X���j��e*�\?".2�h��I����#�Nʦm�{�8����MC��?���?ф��<�V��l���B�O�y4����h�(�D�O�E�9O��O�]0X6M\�C�б!&��`s@��Ϳ�&�'`b6��Of���O���L�A�ީ���]�S��(be�$,�-�i�h|�c�'��';�Ӕ$�����dh�O݋Bw�Wϒ]<�$��bM�M+���?y���?�5�x��'���O�t%�z9�����,-?ֵ��iD�'�R��'�^�8�'�'�2
64��k���<f&�S����7M�O���D��ǟ���c�i�� �#Ί-���zCZ�k:��tk�>�Я=�?�'nA�<���?i����=���`�K��e(Ύ���7Mu����p��Z���t�I:-b�0�݊��"V"ݷg�Th�t����T�w�d���4���9�2MP@/�.|&�0�7�֝y攤)vS���I䟈'���	������<�'S�:�C��GD.�@[a��A���<����?��f+�O�(�'�?���ȕ�܀�#莽;�rY�+	:v&���'m�'���'�*R�'-�Z�2@�,�"�9�"RaT�9l�����I�������������Ov���*X<��Dl33s1j�c�H�%������Rсg�$$����C|0�i�8F@ա*�/x�BMm�y����韜��4�?	���?9��o���6"��q��*Ir`��e(�v6M�O���ֆ4����9��|�A�����B՟h�f5QAa��!��(Mg�2������@�I֟��M<�'�X8Bң��\Ƥ�+�C�|���h1S���	m��|��M��<��2=Z�"#���,�Ā#DA^`�H�xe�i{�'��'W*ꓬ�$�O��	�>㦄X�� '���@�"�(n��7��O^˓q|f����Qͧ�?A��?7��?p� X�3�,f�ڱC��M�1ڛ�'BC�>A+O���<I��CU�ϰx;�K�d/(iF=���K}�)�y����r�'"�'����u��z����'�ΫD�>�p0����MCf_���'�]���	̟����B�81*C��9�S@I! ��q��w�ʃD����I̟L�I�?=�O�2�S�jn�̠a閩8ڔS�'��^?�6ͬ<������O.��O���;O�x6��>Z�R-�V�W�(�|��P����O(�$�O�h%>]�����>f�4��SG�NlH����M�¤n�ޟ��'��'z��V��y[>7��ǖ���n�9Rf"x"��d9�&�'��%���y�'ƈ�'�?��?�qLJ�Y�ޑ��@���m[VL�+�I柰���p25!a�t��yB՟�y���|����0+E�r�dH#��i#�,:�')bw���d�O���&���>��4�@�5iwUD�r��8<�0n�՟��	�T��������OB�'Ds,5�;	��`���f�*�Z�	�:΂@nܟ`�I��L�Iҟ@��@'?���H�y�D����^�.l(��G8��� Hh���!������g$/+��b5؇vjԠ�ҁ�M����?����?��x��'4��OpL��[9�sGbģ6"�H���'r#|������Iӟ���̚�v�$�eE!?ke*�7�MK���?�ӗx��'�|Zc�r0g,ƴ,i��B��҉h�r�}�ͅ�y��'���'&�c�� �m0�b�% D�wOn�n��ē�?������?��&p0�F�U�?�ܱ��F̲z����-�<4$��<A��?1���'~���)c��j��A\4��£�+;)�	ڟ���S�Iڟ��	"%+h�h�:00b��_?,�1%-�D��t{2OJ��Op���Ⱥ�(�(�'�?���_�y�,(
H.M�8�bS�$���'U�'H�Y����:���ZZ��S*G�|2%kWa�w����'.r ��y�']*�'�?I���?)ea��o���e�W�r(������fQ���'^�)�ɟ���?7��=NC�y �B��~ �ѭŢa��&�W�pEB�'"�'gb�'Q�����͆;^) ��$$]�SN0�M������"��ӏ=""7Mǰ��X�PΙ,��ZAǭ��V�'��7m�O���OJ�DEy�̟�� y�a&��CԶ�P�a)X� dҷiXl	
��?U
Gek��	3�¤��e�Pr��;��o+��:�4�?	��?��!d�O��$����QB^�d,#vD�j@(�b�5�I*Rl扶2��������؟�Є�I1|��|�7�G�mӒ��q�۳�M3���?���xB�'��|Zc1r�iV-�L�x08�)��9:�{�Or�p�2O�i3&6ON�$�O���%�tc�3��=rF�ST�"	r�)��MT�d�O"�O�D�O�L�J��_4&h[��"��x�#�	q��]	z����O����O$�ɤ|z�O���ǒ#v���S
D t�HIش�?Y���?�K>Q���=%��F$� Ċ�c�09T`t��IE�K���㟔�	ҟl@K|RW?i�	��0����:8����= ۴�?����$�<�tO��O��@K��<nm����R�*��i3��'f
��&�'��Q>��I̟���Z���RD��3����w.+���ē�?9*O��ّ�i��WǑ�;*Ѡ2��?�� �"�z��|)����#4Q[N�g4�x �
ʜt`I����+Ԭ�؇!�f����уN>%����7H�!35"���޶&I 4�ьW�O��I���+%+�=�R�E(	��Z�J�+'r`�s�ٸ:qp c�C �<)�ER F���N	��|Ѳ�JjL��u��1�����'ߨ1JdGW
R3�|p K+�DDzFɍ�m)lAy7χ�o��r�Y�m����W@�m�h'M�7���ʊ�q�9�͂�{�l	�H7@�Z��E�E?�s'��C�R�΂(kF�)�!����4�?���?�,Or�d�O20��ꜧ����GHԝW��	q��ʟ8���F�L��Ex�,ƈ&n��	�m�|h�e�S�%\d�wf޹5� ���s��Q#!C�!CGv	R+�?�=�rj'%ҽ�4"˟]D�ja�N?1��U�$�	G�'��BR�J��?%h6�#��:�B�I�� ��9,���S�
jP�K���?�'F�xC�rӸ\�D��
tUZ�P�hP�i������O��$�O&˓�?I�����W� ��/H�$Y�֪Y$T����+�%	���g��/Z��y��͸=�$���۽{� �qS��`a���ʫ$$��g �xx�����O@�Dō6�,)�D�[N:�:�gZ�*�6�=����V��T�*UH�"0 �!��V�!���ك�׬bvLi7cW�\��$AB}2R�XCe�����O˧˚�x�	p�|���h��h��?����?�ph�,*�F��\�H���S�d[�X�*dM�+���#�A��(O�H����K��|Bv� f�'%�C���ac�]����C���Fyª��?����Ox�1��s̐�+/D�L���X�'O���U������!�6�DL�:�0>YC�x��W,k4���%�KG x	�`���y�&�aӼ듕?�L~����?��� �����՚�#�� �y����0��&,2���b��S����'�"��IΙ۴U�ecAZ0h�0���&�1kڌqԧ���ن"X�˄ˑ���	K�F�(>�a(��'�"�����O؁�2G,��Ĩ� E�z�J3"Of�r���B�IГ@�%��l���*�HO�S�|%�L�F�N�o������J����Pr%�!�Ms��?�����O`�D@7O���0��Z���Bm^���E���}��\V5�T��o�[L���~�N\���>���l�pFS8��9�)Dv?�%������	�Z2T�@�C$:n��R$/
jrC�	!^ Pb�#�����G�n^V����]0�I޴(1\<�3$ ���͠ ��vYZ�����?����d�O���k>A�$�O���%VP��ԬӔQF�تD�ƪQ��|O���d��[́�R
(��IV��|��'�?y��q�0a[�ΝA�<-f��&{�L0�ȓ Ѕ�̔":*�]�� EbD�\�ȓ_�:�� ޤ�{_��(�F��<Y����&�Rxm������|�� ��(`fD�un
�$�yR�'KB�'Y�8�'�*�O�S�)rL�ؖ�T�䁢@%O�Q�l�<��+ۡR�Da���w��t0��JsII`�Fz�Q��gH�O0�$�O�Ĩ|:d˂���h�N�I,�MA��5�?	���9O�P�Ģ˜<{�}���X(��'H�O`Xu��
_U� ��B֥; 2�
a9O�� DM���	ݟ�'?��	ڟ@��%9��asD@%��{tKS�fp������ �<��O����=8~�8ye�ċ*n��q�J�Y�#<E���E\��J� ΉuJ��֫�I2�X��ί�?i�y���'���1e�,�����̆w��Q��'H��&I�<_ꨁ4�E�m�x��������	�S]V 1I׼Pr��l�|�����O��C����i��џ,��Sy��y�C�W���Jk,@z��k%�Ġ�~!Y!��>� �y�T����`a�:{�pLj��OnÄ�'��	�Ȱ+�
���#X�D��!I�'C�]�����=Y�p@����@ F&:d�@)��<�d�3E� =#���=p�Q��ϑ<3Y��"|:��ļM'�����o�=yB��o��pR�O��E��'��^����4Χ�a�I��xAVʕ q�ʩ��^�;�2!3dO5�O`��Z�����F(}x@u���[�0Ų�a6�O����',rv]���@�e��%�����yrm\

��Y�0���VYB|�aD���y�o�
d�\16EȊJ�6�z S��y��5�	��dz�4�?!���#	BP=�' U*ixdS���m��d�OD���O�ԢU)�ODc�ʧ#��l���	w:4��`��Q��<Dy�(����Dݡ@J�*dQ@9hG���x�y�c�I8L�D ڧ	�Ą�%nR�Y��
���5�\���@�#	�`:&H��ΊLu��	��ē�pJ�$ޢk���D��z��$ϓ>�j���?I��䧈?����?92�U�wF q�)���Hɺ��C�+���i��瘧��	[d�B�$��H���P��s�n����2�ͯ*�ְR��οl�j��d,��C�����'Jb�'�R��O<`�ŏ�J�>���ţ��<x"2O��d!�O���U�a�lAѴ�=y�0�B����HO�i�O��C��3��@���q���BR��O^�DN�b�=o���@������'���'mA�W�0n�B�cMS	���q�'#V��W-�;_�a{"˪�n�FM	'��L�����~B��/#
0(��'�  ���*��+D�>o�M��'
����'$����,On�Ĳ<)`"�>��k�ʰ�씘���s�<ɒ��3,�$L	�넫+k�m�P�S����'��/Yb� l�;$�b�Q%l�.��!����;����֟�	FyB�'QB2�$���'���+m�
Xh�I��h����@S/�p>)��[y��C9Ko��c����.=0��p>����8�I�ᐬYG��/8l��N"N�fB䉇	��D�Ѧ��=�0�F � h^B�I?B��2 ��o6�M W�����	���'j�ER��
��O(ʧ`>� ��*�<ī0ɦ=�l�̓�?����?Y�/˒�?��y*�T�!E\v¹���S�R���+���.��*t�YV�0�����j��D:f-�X�'�J�	���h�>!�%�'Z���1��&ib@� �"Od�x�.�:
3���e�*`��L8��'��O�da1`��RU1���>p�8u 5O���Bզ�����$?��I䟸�	 %�4�cU�B��Xa��+,~LAJ H]����<��O��cx�bX�S���f���*L�	�"<E��M\�$���3LB�!�W0\����N��?a����O>����� CVLO�A*dQ��[g��$�O������G��	2��$,)i��϶W�"���?U��ˁr ��ÖS�ACJ�򥉝؟��Iu!t��4�?I��?�*ON�d�OT ��M7Ӑ�ѡ�@�g�t8���O4����'��J��Mz6�C	�Q�՚�'(���a��(�NH�3�-�5�H�P�0Y�vFr��	o��̰ӫ݇&�@hCm��U%<���1D�0vg�A!8�{�-�4]���獐��HO?�	�L�좠I_�Jj�5��*;��B䉼\G�p�OؓJyF�1��:6\lC�I���Cn��j2HA�ET&M`C�I�2�ƀ����W�(!J�l�Q�LC�I��V}�'*ʹ9�R��wHM��,C��02���O��X�p�3DM'8�`C�	�v����4�إ�0�QP(';�VC�		 �`d	�".Ӄ��O+�B�	C�����;b�┓S��rB�	�c�f�����nZd��5��2B��B��&^F�kE-#8�[�#I(j� B���`��5�ŵ%���h� R�L� B�3yxԁB�!FБ�DR�g��B䉬0g�� ���)Q�A�ae�f�C�)� ޭpb臕'�j�*��	��j�"O8���d�S�R@�F� xH�Q"O�4�u�Z�2�,�[ O�[%�5"�"O��
��ů$)��p��G�m �c�"O&����I-f�
��������"�"Oj��.�H���"��^%(n<u�"O8��� �3@�P�9x]~�C�*O:��V��>k։���� K�)�	�'�<��F%�l�,��tn��~�	�'�
��&B�r��C��>�j�;	�'�M(�g�>#0��a&�\�0	�D;	�'%��H`�ͧLL�2�Y;�D���'�h��a�nzQb��-�����'�P	�ѯR�&��.U*����';\\s�,ڹ1��!����=(�Lj�'j�h����6Q�h�B��/ ���
�'�ޱ0C�a���"@ �G]�*
�'������^�h���ųA��]y	�'<��Ê6�`$s��A�f�8	�'	2�k�-Gyl��H��;�d�"	�'G a���NG��E��C����'^��x�H�y��W�ȇ)���x�'x&�i�)�9W����S�!4�4��'���X�oE�9� pZ%!O�l7$�X�'D�ђ��=U��D�_���)�'� DY��^��qY��ҎL��4��'���JS�˴[���*w��2H),T�	�'C塜	W�ش�&�	�0h����'�-;ң�((@��8�F_9Q�Bx	�'q�CgB�j�"��5k�8�6�'m���Vp��I)�>Ӽ�	�'D�(A�n��q���h�n��	�'D�tk ��"���T���v=��r
�'F�Z�a͙�6u�TD�p����'Sv�í��0����3`�7kp�D@�'��T��-c���I�U�f�\		�'&@�`P����,9�NBh�,*�'���󠄤HVr��Cb�����'�(���՟U%��7cXY���'j:��!H�8"�آ7�Q�Dz�C�'5��p�$�!w��%�����ߓb ��OB��
E�Z���gH�1�NPk�"O&ER����?H����[�e���J��X�����X,2��0c2��i����"O����όQ���Z�Ô�4�c�ݭL��O��}�sPҨ��F�	`6E��(!r�:���x,�C#� *�d�a��M�B��I30:�!����H!�5W��+: Q�
�S](���Q���Z����P�Ȳa!T|�Ѩ� ���ȓ�h4�R
�	^r���XN�pU�?�B���~R�)򱟪{�F� ����ь1D0��V"O��ۆ�ȍi��L"4IV�d
��H�i �D�d�����DZ.P�4X	E�� y��I���D�!�ٌk[������.W��j�U��1O�h�E��p<5���K6�����+B�M`��b<1�����2Q%��bq��uf?Wn�X��&,�X���($�~��NAԍ��/'OF �c����'�\��AkgK&��Iμoi��'�>�3���]Vɉ���%i$���O���A����v�2��
!�䙕����"O.� 1 H�zL���O�,E5�<�g�D���Ћ����r���)\ۨ�����y�&��*[&% !���	[�@���DTL���;Q>b�Z����'��=���I�(����\;N�tB�c?}AR�<�,E�B�(����L={��u@�k��� �4��KJir%�O�	s���J�N^�|7�e��.G�/q��2�f�Tn�4D~�隀p��(�~�PK��H�>�z��2L@��c	�t}�5��Sn.:��q�'�6`�������Ġl�'l�*�g{*8X�����oɄq��d�V�2(f��4��ܟLc�]��� ��v~ʟ�@3%p�%r��%�
�d/)>��l9�OH�D,� K�zS�:e%�0����ʅ�rbIsg�'?ʄ�v�'爡QR�P/S����O�
����\�ϒ% �$�r׊�T�\8�=iAM
1��4b��'=, � ��[�I5��d*U.[�jY�Yp�V2�R�dY�e�����Q�Elt#�#U?wQ�<v���9E�\P�N�-�Y��%ؓ!W�H�W��%5��v�ex����_�,����-!w��sN� м��A�'�F��Ƨ�����ef��q.:���1�:���dĺ/�x�;�h�:�6p����0tDy�
�=�8�B��V8z"<x����!Tx�Эܔ�R7���KQ�uG{�$D"u)3���x ��(b�B4�~bS#�8P�B��
��PRf]'��'���[Ӂ�)0m�D��*%*i�N<I��H�!�Y8a�R��:&����v銥S&θr$M��#�XI��8�]*�@1��c��T:����Z(ӡ�43�(!8��_�ɚ��ɍy�`%�#s�60���B�-��ܚ�FP��~���88jP`���35)T7��>11!D1�n�����3�tiP�L��yߔ��P�N:�0=Q�Fܜ/JJP*w/��]t���J1 �t�j�dޛT΄u� ̖b�'
��PEP]2$��.�!2��'mD�R��0_�`�3�� �BС�y��"B!Bѣ�ND�iX�1��'�� �Ƅ��2�AB�T 6_^<S��)̨)Z$��0d�H`���e*�D}2�^N���V�c��u��d,��$�	ߡ�j�8�O�?��y�q�\0��gפV.�T�G!7�pL�S���Kt�ڹt���F/�j`���o[_X��Q��ϖ~	NP��ѲFƾ��g�C������x��̱�)� ���Gg�`�����Ћ3��<�&ǜ
>�dbm8ړ!��:��\�uO��3����zY�Y��J#���r%D&V��ybNI5a�(�$��{fFY!(��
�/n�BePeM.?�Ua2[Y~�0�,|�SG��.'�L����A�����O�5���pfĄ��~�G}R����lY��4+MV�rnQ�<I�&شq �M��lEY~�)M�m����b矪JG�y�g	2*�D!�����k����p�'Yq�W ��9��Q�eLˇgFuȓ� ��?����O:��)�5���� ք�#!��4+�PZq$=�Ox�[u�èga����ukf��U��ZYj��`%�Tp�'4��J%��O�ၤfݬW7
����b�K�'�E(;_�Ѹ�̙w��yӎ�$/R�<��
(L��M�u+��so������˚�����ʁ(�S��'8�hT(�;z+���G�%Ȉ���䗍,/��JP�J)�leeg��	^~�����D����&�F�&X���������xժD�c�m��j_�|��#��-J�:
�Ӽ�Q�� )"%X`��`�\d�R���<�&��OhJ>%>��ƭ������N�G\:�qL�F���yv��2��B���9���0��x��C�QG$�c���'�-Q��~���r���?r�LؒtnҊPiJqP�A_
���̄U!���/ �Ji{T���RJ�!�ō��B��B������h(��
T8j���@�Jh��|��ɠ���%�%lՆ\A���
)�R� ��x�I\yר�΋6n�J�	�"��0�����VQl��.��<9cM��ą�'�L��'Kh�����l�~�(��'x�����h�n�*���4J��p�E�%ډ�#�ߏJ���.��Yp�'b��@��$Pq����U�>��L��z�ܑ{ዕ���IE�v���-	��4mLdh����W>X�8�b̰i���28T$�0��o�q%�#:���*�K5?! �Z���ϻ+J0#�!V�|Kv�+��k1�b�bD���ٙ$_P �F�ߛR�J��?}C�X��ٖG! �FՠR�V�
�N,)���zH<Ѷ�Z.^�͹uB75��"S
S�Ġѩ̾o�I�x��}�'��h�����~�V=K��X�7 0;8hh�ĭ�9�"��2?0xH�D��y9"ԱXƲ���H��aGJ<#�C�PFh��Q�$Vc4��*��Ė��9V�	���'D<��ƋG��P�x��W�O���A�y�V�K���B��+<x�8�U�W)z��`@Y:�yraKQ�4�c" �$Ch�a픁���QCf�`I0���!\V�y&�9���f��>ᬤ�m��~�d�}�
c-Š,C���œ<�hO61��+�\�P�4.#i��M��c#4��r�)C��:�� iZx��	w; �0����<���5���J��K6h/�J�2a��ࣇ�( ��Գ�T!�Z�r�eK�(�J��@cd֗F��A��[������ K:��QX@
0�'���7HB�+��I�0�"lXi�Ó��\�D�A�`1�BK�F����1q0V���@�|��&m�)*N�k�?[Pu�c���<����m�0H��T+u�a�5�b~r����ôc��@�R��&	�I[�DY[�l�1qJ��H��Hb�@��&{!�� �0�E�։O��Y	7�F*H�2� M!]|z������03n�Şd�'̒�c��/8��t2@�I�{E�y�'y�a��C&�pU˰����8v��<!�	V�s�ڵ��!�<���Ak���6��$m�m�#�C�az�2O���g�c?� �l����h�/�fb6�l�<Ѳ��'V�QYgA]&�l�QZS�'ɰ�2��L�O�QSo�%F.�yU-A�E}<�
�'�V�KTb8S|�#�D���R�l��@-v�s�'8�g�B�g�I&l �����-殨�A	N0 �BB�	4j�ap�D�?z��VQ�}d"��7�c@��!'K��p>y'!́�^;��\<*�j��e�j�ڻ|\��$��:���O�6--?���
tI5C
�.(�����N�!�DS�ސ� �9L� m!�aǉg��w��!��̟Hju��4�U�/��ϧ7�X,p"���>��yR˄(JB���~$��ɏ��`qr�
�4���ߏ�M0��X���M�d��L<!W�B. 伳��V%0ޜۖ��Q8���s��_1OR7�F�`�L�����A�%CQ� D�H���-.�VтG�ٱ����dm �	�g���>�~�T��4g�`���2�n� ��@�<�0��A��@�U��0z�����Od�<�a��	6Tqx0,\)z�4(b�__�<�FjK�r)��8 aJ"N�0�сWZ�<�����S�$�R���0��E�7Cq�<�G^<D"�TLE�G�Y�D�V�<�&�I�!��t�!��?ipUB�#�O�<)�Ŋ>�8�H1&�)�.��U�e�<���I�N4��#sCf,���h�`�<��e�����M��P�I���C�<QA�.xɄ��b���"�R�d�<a7���:��YV~�eY��f�<���rg�p�uդ'�4�hb��y�<ApQQ�I��k��6�p�<9�I��QRt�#��I�؈�D+�o�<���u��hT��#M�P	��q�<y�ƨ]�}���Qs�#�w�<���q�R-b�%S�|��lw��^�<�a�4^�h�@4ٱM�-U�T�<9Ԃ�/��MS�bP�Un�DA�J�<1��4,��5C��J�x����M�<� MD�S��M˒�9X��9�'�CF�< �ĕ
zΝP"��z�漀׋�i�<�VJK;:�(p�E��;�����L�@�<QD�X�'4��A2L�Q���3�&GS�<��ĉ>p5
7`>6��9㥆w�<���Ht���8�*1��ؤ�i�<�X�z]F4qaHӫ�6���JRl�<Q�/M���(`��i���[_�<�5�6�>��b�{�J��"o�a�<Ԯ/��Q���o;b4�\�<)dF�l�X��e�l�����[�<s�L�oN�]Q%�C+,�*��_�<ySn�q�\���[&��$�[�<i��/�PK�!Kl����K�<�l��RJBq$ȀIGj��I�C�<a� �l��B�"��A���1�k�<�G��1���Bw�i)t\�bʅe�<��-�t�10HLN�ޜ$�F[�<QS�.lͺP��l�a�|S�}�<�eK�+؈�h�l�m��IP�k�@�<Tb�,}�$j�B�/>����oGs�<�� �0��[0e�!� $�g�<�6��<J8�ki�YX����d�<Q���DK晠`J�(r8��V��i�<Ya��c5pՈ aЏj	֙���e�<� �!�F���\�����C�"O��"��Pc4c�+*m |�P�"O��c����,~��%��u`�3"O���pB�|���Qt��%� �pe"O�TQ§Ɯ\Jn�;���-�^��"O�u)A�9g����9`g���"O���T��7 �Lm���T�>�ƥ�"Ov��@dْ)�(uKf,E�<��;�"O��d�T�Z��P9F+D�"w���"OHq�&��}���J��Dmha�"Ol���O��!0������rh�M��"O�`���U'�4 �ȝ*V���"Ox�W��%�lq�6ʜJ?��;�"Oz��]%T��z&	��2��{r"Ol�V��?
�4�#�_��f�2"O.� '�)1 $��F�<[ŃU"O�D���l�)C�4k�9�H	��y�)nD��۷���2J=�T�ʠ�y�G�"K��P��N
~	$��S�y�R	pd�p���G�}E�$c�-�y�*_i��@zwgɇD�`i#�/�y�$T�M�UY!�;AB(p2��/�y�ϑjT Ӫ��,�`���yBH�7�NԢ���T��!H�yrmU�pkRҔ�P���$D�9�yBg�0xIP��Ղ�w���B�?�y�m��?ȍ�n� ^�5"$L#�y�+�H��Q���{:�8�v����y�I[b�֪	#s����A	�y"$�`�L��7(��d��|��K]�y�R�Y,����C H��腕�yB臕/jȝXGHB���(��я�yR҂@�9�)�w�����Α�y(Y�z^��P�_>o�*lA��E��yRI�MKzy`'eߢa���
熇��y�[�o.�BRN��t	5J� �y��<�\�y�!
� � @@D'�<�y"�Ԯ~��Q�T�P�~��q��i4�yr�[�&c8ua�-�5u�DX�W-�yr�����r������@]��y"��8%��x�M	h�hbE@��y�!Ww� h,U��÷���yB���P����gg��|����ح�y�Fߧeʕ#��� _�:���^��yBE�A�Ή[�BΜC�Ju
�g��y�(�;&c�q�hA�4�
*h6,{�'ׂp���M�$�"L��Kl��h�"O}�۟r;�����ʠk!\12�"O�-�L
�� D
�U��as"O�(�Q��*V$C����Y3����"OX��e�6��P �N�Ȕ��"O�m�K�"��e���M�W�1�r"O�I��L��7Ϧ�;�@��~}�	"O��;�i�,ꜘX���:DȾ\�"O�ݙgΞB�y��\�:R�;W"O�8��
}�dY���i��h�"O�h�à>ӠÇ��3�z��"O�M�ƌ]*EO����#���Ҧ"O��WBS�}��T!	>��@"O8�$�"h��X����"����"O�I��p���Ud�<CO��3�"O�1��L){�H��`�ѷI�*�ڦ"OL���"��=��Jʻ��� �"On�	���Y��)�a�ײ&�|�#"O� �]
o��a$��r�̤Z}h�[Q"O�a�EJ1u����̽f�����"O�%0+��]�F`�j(�z�"OX-ru�/)��ST�X�NĦ�k�"O� �S4RZ%Wd~�~M�"O�S��V;(�v`��e����d2�S�|�C�F7��e�AL��XǂB䉧��pa���0}�� ��eV�aobB䉵t����R�C<�� ��;�B�	�M�����Ņ]%�<��aE�x����>٦哗P�X,�e�?�`%@b��p=���ט^�����菔��)X���b�<y�#L;Xbfb%�:紬�B.�^�<9���(\�+�"|JDKs�c�<9�*����]��!u,�R�(�X�<a�b$}�Y���H6*TI�`��P�<��cȎh5N�C#з[4�( � Q�<�"�{i����eܜ-�r ���.T�P���(�80q�K�0)����`3D��)�E4-�85�7��C�����H.D�,��!_F�XPK�4����.,D��!���)n��0�w�N�l܂���>D����N�g 2t��-�;+\T�sP�:D�,���G'�`9
��B��U���yRo)5�0�!�fR�}�XI�,��y2$��n}ȓ�8sM��z���y�D��4�y6e�g
����h<�yro¾t� Dz0
E�W�zȺ2-��yRǇ2(�t=Ѱ�@��In̰S�!�䃽4�tT��m�Fzq"	E!�X� <�����C1uP
삦�ݘ!��P�%^�I#Iٸ_C~�p��ܞ�!򤕔��Vk��r1&���̳w�!��9�1weWl%(K�m��S�!�D�=f��,9%�{����Ս�8u|��/�O�z�lA������I@��:Q"O�l�#Ɇ'*	9�Bk��%���"O0܁2�O}c���i� \k�@�"O�$�I�4c^�c��!s�A��"O����ΣBQ���6S�UƐA�"O��U��^�,e����):O��`c"O�� �H�jf~���BՌJ��	�"Oґ��P���!��k�����C"ON��cA�L�a�ȁ�0�5�"O2��P'R/V��{���&"��t"O1�%�R�.V��)�G�w䰋��	\����Z�:��Xȱ��3}:Re醯Kq�!�$��@<BP/ǣ|��p�O�m!򤝇O�x�8b�f�A����7Ac!�ė�W���I�Rc�r���G=!�D�J +�gŌ!!���%a������Q̓�d1開��T���s� �zA͇ȓB@&�`��<`� h�� #M�4��ȓB�!��
;���s&B��>��ȓLj�@���Q�<AQC�ZH⠆ȓ����/�iDb��r��C$���38[��<j�ldP�GF�x5��}T|�#�M�:F-���тWڴt��IA~"	��c�ψD
ƍQ�ޏAu�C�4q����	+c��4jU��	!�C�	��~�9r���p���(Q����C�InD��$�E�4Y�x��GR�;i�b���'��~'$�{n��gǙ.�*x��Ga�<�M%&�t)�ؽM��hk�e]�<� �t��BY��(7��.f�l4��"OzU�q�6�vyI�i6P�4"O@ܱ�.�be�#ٲ��"O�D�g�N�9Y�h�w�C�&5Խ��"O����()x�2�i� w<�T��"O�E�0ɕ .��鸕�Ҭ3 ���"O
4�U�R8U�(�s�&l�4Z�"O0 �+̬Ao��ӁU�Z�;"O�hW�P'�|#��$U�։*r"O�j��� x�@,�E��6�n��"O���҃R2��9�MLJ�v ��"O"�!UۗW,C�k�Akȥ��"O����ݔH�"1'�Ϟ1�X�$"OZ����._�&�����7\~x�i�"Oe	0�ȑ�������5�-:��x���[���OX������2�'��A%�4��'X
�r!���i�*m��K2</Hd��҇�HX��b� �06���	� �!7��e���0D������eCQ���qw�ih<ib-A�':�2b�=5|����\�<�A�W٠�l�lF��Q�X�<I���r�(�"�%H�?�����Mi�<����w\���O��H�c�96�!���hV�`��i0,M��͇,�!�̬L������@.����`@ .�!��4}�� kեҾ���Ư�Zm!��t24u��!�P���DL�NZ!���9�!�m��4��%��-!?!�D�d�r����t���X���/3!����/c���Ug�N��������0�!�DT}H�sq( 99�DdA�J�!�D�"v�J� ߏb�1���3�!�D�/��dPƩƉ]���ꂍ�Q�!�NaF��H��G��hA-P�!�d�����#�U�*��P:&�K�"�!�՜\�
L��E٬L|��5�o!��D�����&Ҿ���>=!�dG�}X�t 5%��9`j��K��!�D�,��0�E͂�T���>;!�d�F~!�3��'�h	s�ڋF�!�dI o��ۑ��*3��!��L�?�!򄏲|�8��S����㞣*�!�$�C���U�E}��#��!�SvSVUY!%F�e��x!�k�p�!�$�.xHXQ䋎�w��Jb��=�!�GQP�P��� ��Y�c�ɻz�!�&,l�� �G�]���H<R�!�D�M�H�)[�� �����;z�!�$�}DDU�fkH?��3��P�!�ܐU�����2h�n� "E�!�ςX̸���=	ͤA�7A5!�$L41�X����lk�=�#O,�!���yTA��QUj$&���B!�ٌ]���2��(9��a���7!�ƕk�� �w�B-�J��!���U���j��m��y��
>�!�$�7��%�!h�8 �:�;�n?�!�&*�<��E�3`���0M]�O�!�\l�  *^�b #��!�dC'K���I3N�D�|t�&cY:,!�ׇH�uKM�<ܘ�'(�A�!�\�~F���ԓT|���!}B!�A	�t�bW�E<D���� t/!�ɕE�h�)"��?��lX�Í�/!�� ��i�J��mx@@��L.��"O��Hd�V�"�U<m�1Y�"O4HR��'���[V�f�h7"OrM8��ʶ5X�J�"��y� �U"O���M�+�\�s��!&�0�zg"O���#��s?L{�Z�%r��AV"O�Dc�aOJ;�@�F"`W�=p"Oةr�N���*Q�a���Z!��[6K�`K@o9�4X�<w�!��.u�
��h��Йh����)!�N��C�������ckĜ!�E�g�v��a��b������'H�!��6
�«S� S.$�����!�$6B��d�3PRΰ�H�#f�!�dA�}hL�i��l��aŚ�.�!�dǷR�(TCbc��ce��8�A�11!�$��@&�9a�C�WL�dCF��v�!򄂭w��mH!��_L�2B��T�!�D�`�8Qq'h��d�R����I�!�!�DK5b������6�}�4�ըXb!��$CxX�nӕy����j�;n�!�dH8�.<zҧZ����;��ǎO�!��Q���q��?C�����E2�!�=Di4��LU�-X֥!Vi�9�!����*i���;?��+%��!�!�DȎ2��pA���(u3�u�d���!�D� ��*س2�!��':�!��P=��H���s%xh�2JI7#e!�90��[�-� �u�'̟'&w!���V�q�-��H�1ih!��0dX���垣9꒔H�! �N!�$�	
�:����Y-b�{�E� A!�Ē�5�|r.W�;$ةل�9*!��ٌ;}��2��ҷ#B R7�$�!�!p.���"WB�u;��!W"O���K�E���N��=1
Pa7"O 4떁�^R�Y2��J&+-h���"O6� p�\�(Q&JE�^-$��B"O���c�-O���c�.P.@����"O�E�a�O�c�]�7�N��p�"O���bg߼'�r� sd��BIȴ"OP��2�F{�)*_��YT"O0��cG�R�"�φ$�~�U"O���É�����J
bB�5"Of�1%�؅0��Mk�GS4B�*U�"O����,��M��C�P�Vxxp"OR��3��p�ٲ�$V�9�J%��"Ob�k��9=�X��w� ^0h3�"O\$���+eF�� �KI@�ZC"O�`#��ߵ |d��0��= ��Dj1"OV���J�o�<�s!�$Q��"O�����[�1V�����^X�"O���T��3&���@]�1XI�&"O�%�",��2F�[�J@�rd�lP�"O�#S
��2mn �2j��C�h�"�"O�paW�#Ui���1�G,-\x��"OL�P��5�p���#�`�7"O|�栒�n��P�o�ZL�"OX9�¯�	̰a'ϊ?s����"OT���P���(#Q�B��l#�"O�<�B#a�9��L ��(����u�<y�Gؑ\�@P���)�$]Hp�m�<!rǺL�0���	�M�|�W�e�<���4u9���K��\i��&D�� �ɚP��`�pAC�6
\v�"OL$����(W�@�H��/H�к"O�x���@z~a*�h؋;���a"O\���[d�ЉS��b���"OX$��&GJѡpL�6r��h8�"O�$
���tϪx�)Z�8�q�6"ORt2W)M����2��0."n�Y7"O����;���4��Uz�"OZ��P�?W�:Y0���14c��t"O�Кv,�&~+p\��$C5j��"O�8w*�6�@sĄ�5r1<��B"O����-V�r,0@	<O��I��"OdYc���mf�lIR(��g�<p�"O�%�5^��^�@�I?^�$;�"O�U3�k��)���]�`�Dig"O�i��d �Ll�[� �IxU"O���6��X�(��f�>�2p�"O<����N��W��dw�8�"�d�<Ywar��ʧ �#K��BHOH�<�P�K-K^y" �Ũa�*���`AO�<�@̛+k�������-A��@f$I�<!� �6�MI�e��sPɡ�(@G�<DKD#$Ȧ�	�擀ba�]����Y�<�QJ �:pXg�K�=2h�"&EY�<�0D !$^蜒w��"+CTY����<I2%� M��I�Ԣ,��I��O}�<ykQ=G礡U��,#�x��^v�<���H%v���>1�� d��o�<��'_4O�^���鏂"mL��5�n�<!��$z	��R ��{a��($��U�<�f��<g�&1�@e�
.�`ҕGLG�<��D.'�VXpB��Z�d	C�<�֫�T"śQEҲp�x:u��}�<y1�Ǳ%�2�bI�/yvܐ��k�B�<M�;.l�q�ܦ�Px�GL�t�<�"#B�ƭ-��y`���;� �ȓk($к!����I����"6���S~,�ia� �t14�N�箸��
�`,��ǂ������ H�M��݆� ��gň�^sd�Z��^�%*~0�ȓ>+^M[�J]�)�|�v���U��hNv��%�s�2Lr�~aD��ȓd۔�Q�'4=�<���I5�v ��{.�af�^'j;���@�ش$K�t��,�@�qlPx�R��`�A�>y~A�ȓK�����h�,z����,Z��ͅȓNӾi��h�,o}\Ik�a�?R|���qބ�#�
�j��8�	ѼG�����aj٩���I�a0q��"U��0��f��uP�	�,��$J��A�ȓ;�sE�?v��z��/����'�T���H�"�����V�9�ԭ�ȓ@5�̑��D-���j���n	���ȓ�Z��	#V�r�t�<# ��ȓp�|�S��'0I�0�r͌��Z0��fe��Kp��>[۠����	��x�ȓTǘ��vK��Llvt�5B>D�0:�g�$��P����B�*5i�b:D��򌖼;6�3����*�(��o8D�����*4 �JdN�"E�)8D�����L2Z� ��5��	'���V�5D���F\�<h�K��>m��a��4D��E!H$k�~,SR�L�ba�"�6D�X���|�L
�nK��d�+�l5D�� �Y�IT����Π@&�x:q"O*���H;o�D�Y��� LY��"OƵ1&��6m4��U��'jR(a�"O���=v���o&g"�	q"O숃Qe�$��z�ȓpL@���"O��k�+MWn�S�EM�3VqZ�"O�0��e�>p�.5�FEơ'(`�؄"O����������J�
NF\�A"O�k�G���hx���)^����"Oz*�W2d�V�����X���"OV�Q�KW�-����� �M�~l2"O�%�����$�
�"O��s���q�t�!��F�|�ir"OD��Ǉ�-�	d��5/����"O��0��.���#NG�h;�"O6e�%ʳu��dQ'�C�'��x�f"O2����0D)4,�$��#��M�q"O*LۡHF�x�1��*ҍ1A��3"O4a�`��$t&����
'O0ԈS�"O �j �3b �x�g��*�:�"O��[4��0\l � 	5@hyr�"O���� р�NER� Z��m9t"O<�{0�3���Bp�P�F�Ɲ"�"OP�P����4�B�oi��$"Oh)ك"�+}j�Y��.\`�L�r"O�ig�F�]����aB�Axn0:�"O�����%��]IpAʵ��:��<D�����-\��ó��HI��p�8D��x�!�
O$�(�6��(�`��0�;D��JWj܁<�\���J�6�.�	t":D��{��C�!YR$ǛA��p�6D�h�"c�9���ළ�)@������2D��C�_�p�!
�"®��/D� C��fZ�u�HJ5��(-D�EI&ZN���-�/4ڀ�v1D���&�C1#��jTBG-9kb=J�o0D�+&Hn`&!�0@D?Bf�*C0D���H%z�)�)ys����*D�����E�B�8$Y��A�#��q��%*D��H!i]��m+!��?Yw�-���2D�l��眾#��h�`���J�+$D�h8�f~��.T.������*�!�$ފVv�ո�a��),�o�M�!��
w�T���ЂX��S�K�9�!�$�	�pj�G��Eg��um�[!�dƓC�n�c҃�QI��KR���C�!��ղ?��1S�뇺[����+ƅ	�!�DVX/��d�6D�XmQ#��;l!��'�]��ҝp�p:�'�,,�!�d��6��k2iF�H����FP!�$�2�!P��zk6]���R2%!�W9Rf"ZpO|��'�E��PyrZ�6D\���u���H���y�N��y�F��Ĉ�se@��1��y�.�<N��(�/� n���p$��y�c��t�A�&Pa@1�����ybl۲g����V�_�E�$�����9�y"��i*V@�PC=�i����*�y�E��k豂�W��Ht���y�-	�'W(Y�q�R�&��5��y"AX:_*��Z"�
ĪJ�i���yR�X
�fҁ�ԋw�9X�eM��y"M]:��Y�em,�I;Q����yB�X�I��M��F�=aݞ�� +'�y
� l�ģ�*h�٪%�Q��	��"O. �'쎆 �P���c
�+�px9""O�l�i�#|=�4�[�,:ve�"O�J�OI�+��81���"�D�2"O`�)���Ȱ7�� K7�0�"Ox��孍�>�Y�n�V2�}G"O�@�Jx��e�Ê[L�z�"O���4��yON���K�<&��ځ]� D{��)ǜb�L��0ԭT�Zd�� N/p�!�䖚$�f��掯R���bd��@�!��ܴ{Ш���I� 5��GLT�!�d_/&&��)��j��� ����n+!���d�������G+8E!�Ą$=�6�#�C�N�R��$a�."!�אBl��[�iP��Ȍr�C^�!��K*32.T㰤�yr��Q)�6=�!򤓱KX���M� &PQ��=(�!�>n���@j��Y�48�	�
�!�ʙ�t81�9!{H��'�Q�!�D��h�Kf�
�AB( [Aa�%I�!��SHh�$Y�0;fT�Y�3!��Y�"��lR�,! �5F؜/!�J�l�j��W�.qr��\>6�!�\� �j<TǛ�t����cٞ,q��$�ZI��E�D2[��umM�y��' cV���MJ�5s�؊6�F6�y��҆X���j���64��� 6�۞�y���(�(sFI[�$ܠ�N���x��>>#hC���^���T�I"C��ٟ��?y��D�2�ݫ�f75����F��p�!��՗Q.�y"�oX�F�sgl�!�*^�l`��eR�EL}!��^�}�!�C�Gn��7��<w���͍�"A!��>�NXSu���X��Yp�#D>N!��Tm�fɟº)�#\�A�!�$]*c6�xQF�!TR@��a��{s!�d?N�:� �o5LDp��B�[�!�DP
w	zi���,)3v����<=�!�$"u��Ҫ�m0������~�!��*&���e�;d��R �#'n!�$O:NM��1AKB5`��9p���AY!�X4b��U�p�Y
k��(�o�=<!��ك_K�����">�����-�s#!�䙊��<�D	�4Q��qX��ۍ1{!�ڷg�t�va��FL�U��Ķl�!�G�Uݎt�Hَk��B!�8X#!�d��h�2�f�����P!�D�\���ꐯۘR�\a)tmH�	�!��C�6*`�R�.�����O�!��0��Y�W�J�m��9�R�14h�Oe"�N����)!�S/g�!s�"O���VQ�2�H e�&S ����"O8�6��X���fCRv����"O�T��.G� ��I٥�Z�V���"OV��G��?)F�PkWmݼk�:`"!"O�-�&&M>���vLG@u8UK"O���fW]�4+��G�&a´yQ"O�U��	5-Z�s�N�&O��P�"Oi�R"� l��i��*�U�\q�""O�!B��R�ˆ= 6��#0��Д"O��5*G�L�~���>m� )�"OX@J��V{�M��v���"�"O"4"u��=R���e�bMB��"O���wj����N�&I�DL ��'����i�? �@0U�0ڜTꢍ�D�$�"O:q��mM�VYm�,� C����"O6�y��V.4qf�̸B�N�( "OJ4�eȆ#r�x������HF=A`"O���Ǧqgj�d��;7e{�"O�]�0@�~�Da�te =b4ӆ"O��C��#>te�µ�P�^����0>�P(�F�بCBeJ5�0���F�<тh�))�N��c��U�z�Ey�<� L*zc.�#���&3�Nᙗ�{�<�3��@u�0L˗n��ɶ�|�<IE��C� 
����ag�Hx�<)Bn��E@��R�Y7l\��P�hu�<��� [���fش�DU;QeLt���0=��
�Oؕ���)0Jɫ"+�o�<Aǣ�&�*0�-k��q���u�<���G:ھ ����(U�bD�F�r�<aK�b���j`@E(Z6`H���j�<���]@"F�Y�9
̔�a�c�<1V��o�B��G�q���q!f�[�<Vʞ�"b�L��N, ��9�T�<��b`�)3�$ּpi4������t=!��˧p�:t(pK�^:��p�J:!�K۴�I4��tY�P0&��.#!�W�r��m1 �Vڀ2�`��i!�$ʸ<"�$c'�]�X@. ��	ļP!�d��W��X#�6xty95gZ�|E!�dЄz�p�*�A��#��cd�?:!�Ĝ	g��`0�^2�`���d_�B�!��$/��5��MP�^ˌE��"-!�+/,X`�`�D�����E,!�D�3�L��$,ڢ8��DƘ��!�3ײ�t/���ꠊ$Դz�!���{���-�Dͪ�:2(O=Q���>O���c��บ�j��m�h1"O�q��m����Q��ꀘo��Ł�"O��
�F�?A�(���)�i�N=y�"O�!�� 	PzF��C���	:"O ��W&ޤD�0E37L[8P���0v"O*����/����K��i����"O␡��߷��MAĊ�&\�n1;�"O���ȍ4!$���/rh�H�"O> �P�V�~�<�x1� �0��"O�i:�@ڝ4��!ph�KǬ�ز"O��5E� %d�yn *_�Pd�"O�h1���2��9��Ԥ9��"O�1�bG<;�"�Pb�Δg:��"O0��b���65:��B=�����"O.�CI�y��E������"O����ȈzF�Ap�L��i�X�	u"O!���:!)�s)X.���"O����G�h�a�b;).�-�"O�٧�)n��aJ%t��"O�EX��Nw��	Ɉ4r��e�"O�x3d@�0���Ň]�L�<q����?�S�Iו9^9��_1xҥУOI) g!�D�WD�D��'B��"�b�D	;Fn!��;#��VC��]�0��E��
�!�$�r�	&�Â<���ɧ�Y��!�ą1o*��6�Ӭ-�Jh3�	�Yg!��G�D�����8Q�(�y�n92Q!���+@*
|��F�J��`���[X�O���dy���eM�h@�.�|S!��M�9��`���Аv�� ��	K!�� X���K�?t�@�� ��I*%"Of ���>/�3�A�\�F�J�"O�M٥.L9P�<"�S�ivI�1"O|�����UH�C��T���a�"ON���aCd:  ����Z��	A��{�A�s2�� O�)SmZ͋��=D����I�!��z���\�	ۡM;D�(H!�xJ*t���-�>IђC8D���t���$�V��$�� I(����!D�,�e��,��u{1�ڹT�&B1j D�p)A׀B��tN��}�D�&�#D��H�+�6V����,����n&��4��V�'�:�M'dݔ`k�h�1;�UB	�'�D�qJ��OY�Ӭ�Whi��'`�hR�H\uL�#��=Vx�	P�']�$���;(�I��ɩL֢�`�'Rt�ԯ��8AAhۅH6`i��'����#+�ŉrf�UN>s�'+t���ڛ+
���J��C�@��2[���'�ў�O��������s�
�u��c����'`�2pkí0����	G�BpR�'�V1��/]+k�.mK0�/:h4k
�'?�y+��^8�n��	Q5-�(�	�'C����^=&pu����UyR�S	�'�(
�o�pBҨ2Ԩb��c�'h�8T,��8����W
�,,6@�
�'��|GkA�9����݈P���
�'�ա�IZE,����d
�'mp���� �JǍ��D�P	�'��� �ѧ>��u�Í~R�ݓ�'�xL�G��'g���0��' ��ݘ7���x��˿	ƨ)1�'	b�9Gd���q��!,�*L��'���dغ^Fl��`F������'E�h�����6S� ¤D�4ҘUy
�'�����%�̵��ֱs�2�p�'�A-Ψ3~��ġ��q��:�'�:�b�	�4�C#H�7~Αk�'���	���4ኄ���T<x�y�'���2�
�F��D�s/�
"4�A���yb�D"���OM.7�lpfKܟ�yR�^49�����.}\H)XդE�y�[�*ɠ�Z$@�%����W�yr��:$Ԕ��aN+J@Ը�w��9�y���y
z]ktK_�j�$$yg6�y�
B�ƭ�!F]�b�APG�
�y"`<e��0FK߸F_:����yR �S��
ƀͧT/�0X����y�l�q��ՌۉQ$��
��(�yB���vTz���H�D�H�E���ybI�S*�p�G��=�`Xs�7�y�o5���4"K�:���1,Y<�ybi^�B�����R0f�a$A��y"k�;�X8�A�;~!(�A����y2�^`+z�!��	"v5��ff� �y����������w��Y֪�&�y���Ԡ{��\���Fb��y���#!>`���.�O����֍���y�n�.B"ҭ1��]
4P��a��y�cΊ�R�r�g
�W׈�3��y2�Co0t["�,GL(#���0��=����$��4�u�H32u�ez�$;m!�D��PdZ�f�\�q�夀!S!�� rƀ"��c �P�CD�|"!�� ����P�}Ȣ1�c$�X)$�"O,�h�D�xU,�h�h����x9�"O �	�C��%S#M��LU�d"O�1��� b=&E��?�Ԡ�2"OX0b@�ϵF
q�!M�s	��	T"O�����W�'$���Y��l�Z�"Ol��AG��KPęy%�?о���"O��KEN٭�-Z���b���"OP�Q�DPx��yw�A�PJ�-��"O�,pգ��F�d|��_�S�l 1�"O��*R(���]���ґ9�z|�u�|��'V�D��j���[;J�2b�^�q'!��^��,���Ku����Ă�M!�d$bY�<z�K��q���(�q!�dU�E�v0��*@3&��i��c�!�B2\�-h�I�<?�a�p� -�!�Ĝ�C���B�%����Y�Q�!�$�f��,�$��9&JT%Z6?R�Oz��nG+~n83!�,8��#A"O$�x���6Er�W� �)�"O����v�"cD��k���D"O�i�K3l�����h�B~��"Or�r0K	)H�X�ǘ 6��"O���	ֺN��$B$H̓]��"O�p{�B	5�N=BW�¶2�4h�u�	N>9*�� ��%C���;5�u�@�!D���"��7�!ˢh��(nRl3>D�
�#��%q<)[�n�=t�>��b�:D��i�펷9��	��1A��X�:D�(�w�L�@���Й
�M�SL>D��
dG������d�9;�� ���<D�(���׷q�t˦h�(OvPuM&�����x�%͍�`(���FF�t}
���"Of	�*���Z<� ��4qČ
p"O(�XG2�����Я8���"O8	j1��A�#A�)Gs����"O�dBJ"��ث��E�n5�V"O2���u�05b�e׽�a�w"O&��5�]�Texx䦞�:!RV"O��󄋪7/�QC��� T�FY�e"O�Ce��
^�x�a䋲u�*(�F"O�hR�-��Cr��tL��`=DQX�"O0h����"�R�hU.A.w:P�#"OuI��a|��{D핒ET�)"OLm�n��ZV>a�C�8n�풗"O���*�Qv򔣀-I�K�� "O�����ܯq���ؒ��-.�X)qV"O���  ��SK2�U�y�r�"O`Iq��6w.x� �U	D�2�:b"O���j��V���ӂ�S�t��"OL�� ҙD]$m�g� �hD�p"Od����eJY��FH�z{��1O���T���s���c�B��]C��O8�=E�t7O,U���U�<�"eK��	]*ЛD"OL��3+92M��[D��5pP�l�$"O@�xr�TR�w�,'X�AE"O�Dy�!ڛX���qi�]�&��&"O2�hG��+*Y��
L*F�<�B"O|�f�хx�6��%��.vVP��"O��À@��f�tU�ehI7p������F>�5�<`����W�M?8�&IW9D�B�%	����£���EId(�e�2D�Wd �/Sت�D�:a���0D���V��0*U��nM�"V��*<D�� &�k�O~ch��Ԥ	���L�"O,ٻC��G���0�+�&�3�"O�i��[G�ZA��"�7��P���'U�O�}�EKDpc�%�Q��C��!>l*,��L���0���*6�y+&$�2+L��ȓY,�P�* 抬�􄇗&�����8Ҥ��d��Ij&t��?s��Q��EL��6�1(��t�5��c�l �ȓ;/� ���\@�=p��+8ߚ���Q� i��-I�Qƚ����(#�x؇ȓ6b�x��J�@I���g������<(�祚�
^.TaR`�6D����UST��F�O�&[��6���0ݘ���u�ބ+���-Am�
V(K� �[�����̀�h�;�L+�d�ȓ6�z�aA��-O!�Q�ȓ+����t��b`�X� ���i��	� �B�5sf�&�ŎU�fh�ȓx ����;۠��*��[��U��9���cx<4%��K�\0��(؀�H�ǔ$*d5
�郝V�̉�ȓW�F�z��[ pEd��/QkH�t��(�d�gdV?0���p/_-=Ld��Sz��Q�N�,������$��?y���~��bj�,t
�挲[ �Ѱ�/�K�<�1'Ю4��<�,R+!~����~�<�৉57��D�w�K(8������W~�<A��;!؈I�v)��LS2�ð@`�<���� $�Q�E�o��u+�`�^�<!w�O�r�68hu��(�R|�sD\U�<��o�'r���!�jˡ8��e�&��H�{y��O���Y5[R�B��Uw<��'����Ś?�.�� ���&�,*�'l2�9s�<z�A0�	���j�'.p`bn�B��ь	�� m��'������ǥ"n���M��	�'��A!D�@.& 0͞=n�6�	�'�dh�A��T(dKϬ;�(�L>q���?q�'DZ�����V��ة���x{ָ�ȓb�0@�í��9�� `6Ĕ�> ���z̫��L�Ov�=��o?1Z��E{��O�����ŵ���;�h�v#��#�'���a�GU��`�Ri�w
���	�'�T;�D˄&ܢl�R��&z����	�'a���G��6W@H	CF��P���'��d��:4N$�����w��Y��'7��0���-(le��_�qZ�'� X3�֦a�����d��^�"���r�)�T�����Y�Z>��� ����y��Ʒtl���G^��9��Y�y�C��t�r=
g�T8j`������y���J;�ٻ���6�Xl� ���yB��;b���J�R42_�]0���:�y��2��<)�a>3�F�KW�	��y2$J&A�@pC��3�hu"� ��yR��#L����^'d�հ�װ�y2f�4*,P	)�a=$���y��^�y"dɱdd���'P@�6#�yҤ��Q*���冎�}�(QHW��yb�"_e� ���,ec
��3�yR䀫|Q��P2�ݎP�vx��V>�yȍ4�����JZ`����N�y"kQ#P�b�ç�J�C�z�8�c�<�y�×�	:�<r���r�Z!郬���y
� f�WB=����&nٔLT���"O�9 ��[�n�8T*���:]�ZE"OLP"�V�Q����M�,ޕ�"O��cL]��&$��A�'(,�8�2"O>�"��I�-jqx�g�9�jQ"O����H	�P�� �@��'r3D�4"O��燘L�E1`L˒Uv���"O����+I�>���r��]h%��"O0�Yg$Y&,@t��ԩ��6`*��"OБ�hT43*���gC�d���f"O<�F3wkН3���c�xă�"OR�aD�ԋ2CdT�U��LtH4"O"�*"#�9�ꀯڅ0b�E["O��X��i�዇.�#([<���"O� ХI�J4��1�1Jh��W"O1�S%�(cUn��I.�L�Q"O4X��T�h9)�\�O��"O��S�ċ3���$�#m�݈�"O|���O��՘�Ň K�`�h�"Oz-��_�q�"��������"ObԹ������׬ؽ+q�h��"O`�x�d�n�^�{�ID�r���s�"O���d�����a��7U-0 x"Ou�a 
�@���G�	#*��"O�0fb��>~�)jf̏pT��D"O���:��3EX5##޽aW�'n��{�j�P�6�1���.�B�|��!�L=��`�FI�K$�B�IT�[��� 3�(�'�G�]i`B�I�82=:�Ƶ6��!AN ��'��'$���q<\������:3��3?�B�	���\9��҆{��p	E�V�!��B�	cz>XZ!D�>gCn4�A,W�-n�C䉝LaC���mĈ=�07o�C�	!� )���̹<�& 2�h�QʢC�*/�fYȁ埅a��-[&�
�HB�I�3*,u�m�
Me�����Ǉw�B�=1ç	�����_�o��P�)ݕ*J��ȓ*�.@��$\�Q��;��]�@yꄅȓd�����׮.����S�Nؼ��l�'�I� ��2E�
u�+�J�
���'��૧-� ��ģT�[�<�%��':b�1B�� 7N�	���R9�0�
�';�]Q��N�����+g
���'��=���h���1M<f>������-�Of2%d�[��Eb0�&?�L��1"O(�it�y4�-��(N)lA$8"�'��ւVC �\�C���vر�L0D�LC�� )};6ahf��<�2�g1D���"��^��;S�JO�H��V&$D���c�X?K�#F��@��2�#D��hTE����;��B~ }z�D#D��[��_�1�����^8����"D�Ljt�
b���rK�|[8�)B�;��8�O ���jJ�k���S��W� ���Q�'��'�az"3��ESԯ�1S�R�@w���y�o<>fʡS����)�V@J��y2�Z`B�Z�mZ��rh��"���y�ė&n>�E��$bZ��%녅��x"�>|.�eçA�}FpY0d� ?�!���&�	S�.).�@+Xn��2?O�Yɑ E�/*��8`�է<{�Ԃ�"O�4ò[u�d�G�.jd��(v"O�\�tM��h�NI � �+��XJV"O� ^���Y�L'
ͦ[\(@9q�'Wў"~
�&��c��qJAf�]��`����>��O��L��}�RA�D�B���R��'�1O��qSaN�U6�)���l�>�""OҌ��߲�`YjM�Y�@ A�"OT����"R��y�C�:q
H¢"O��g�<@���l� \ ���"O~��U	Ҫ ����ȲD�<Br"O�1����h��!S��V�@�;�O<�hb�:�X�Jc�B!#�a���)D�؋EbL�_���#�J� D�81X���Ov�=E�4� ��@ȓ"��g���1�#[�ўD���),�� �@�,V4 a iB�I7P0�(�%�� )BXYb�Nrc�C�ɤ\Ƕ���bK�Y?$��0��\|B�	48Ȓ$&�"��ӆ��H�^�O��=�}z��5D~1����zL,R#!�c����<�S�Q&H�b�J��<�Py�v�@Z�<��.�U����Ƿ[�t|��PA�<����^xd��Ǯ Ը�Lz�<I@��s���۰	ݾ[�N��s��o�<і��;�v4��$E]܈�� �i�<��猐U�FU��j�$g?��GQb�y����y� |���D!�7
W�3"A��yB��B4�]�4C�	U���!����y�IO5egXT��)�q�Jx�(���y��
XL��
f�Z$�	�㗗�y҄W3:��;���?��Z�JX1�y��]Vx�+v�!C�2�#�$�.�y2LA���S$��J(��"C
�����?�S�O�B���dӈ���I�'0!r\�K>1�����W�8p��!A5*���+3nD�{�	S�'V�	j~�AD��'��6^��9j�(4��7�O����ʵ@��P��]82��ٶ"ON��rÆ>.��)b�#)��Uу"O,]!��ҧ.�3���:���"O<�;���"4.|�I0B�lNrT�q"O����/���s
��) T���$'LO%`��Ȟ9gnY0�m:(!�q�'Z�	E��!@���02�����Õ*�jB�	~�nT���Q�:"<h�de�3Z��C����)f�U��$�xd��C�I���И���//��*���1+L�O�=�}��e��v=���4N��FH�;EQL�<�F)�̓F�Y��
��a��^�	cy"��<Auh�>kk,!��R:x
z�zĪ�u�<���I(b��z���=�vY I h�<��IL�D�rТ�C� *^�8c��b�<	����F��seh�;n=�U �e�<�1���{��#:%6H��Q�Q^�<���O*;^e4��7f���P�/LW�<�Pn���]��*dJ��fT�'z?���J�3P�4�b���q53A�5D��֭�9@zU�������H0D�Ԛ�Gȗ]X��1H"�V����-D��EB�$9| `r�	dv��+Wf)D�ҰMΙ<���%N�.=ߦ5��&D�����f%*��ϡ
��	y�.)D�KĄ̱)�q�G�Z���%R�'$��s���S1X-RB"W�c�B@8G��:"VxC�I3���r�! 
]z�d�ۆ9�>�=Ókgt(�d['�6�*7	�W?��ȓC2���[X�H`�0��,~g@��[�JA�B�V��%�E�)pw*���S�? ��eN5a��FYp�k"O�╉�3~P�D���<`bMqC"O�`�5bNt:�Ț�j�6R�-�3"O��8���2�$	B�V�.=<Aa�"O��s�����h�	ڪy��"O�ca��?`�$1Q7F+'/b���"OZ�����6>� 1ж���l8k�"O�)��c�V�x�#^�G� ���"O2���
�[P�A�ǌ�c�"O�ܰ�Nޑb�uX� �(��B�"O��AG�L�N�<�h�/�'h��� "OV�y�^�0^h���(ձ4�Ŋ�"O@��s ��&��+���H8�P"On�U	����P��V#�A� "O
���	��J�T9"f���0|�`4"O8ͻ�g^5-���!������X�"ON��� �) ���j�	Z�r%с"ON�@�FJ8.��J�U
q���"O ��p �;HK��t�B `��9�D"O&���=�V�S�G<>��ͺ�"O��Z�)ɋ4%\Idj���Rб"O�a���&i�� �o�z�,PQ�"O���G��gX�L@���J�l �W"O�Eˡ��8D��Q�����ʁ"O`��vO�<HH�m2���w"Olpk����+"��b-J�i54�"O����@��2�j�ړ!�sD"O�1X�Ѫ�A8b��x��""Or�UGؘ_jj��g��⁣R�y���,���7Ǹ;�MAՆ 7�y�i�="�:ӧ5����O���yB"��By�r@T�=M �j7�y���Q�( FgX�-c��:a�֑�y��6PW���)��0�0i�3�y�$D=�a�V��5KXd"ѡ�<�yr�V��\"�]X�(�˵!��y��W��*G�ͦz�VQ�$�șE<!��E-�rŌ��0e;g)Y8B!�$��jM2�G\�K���:q��"3!�$�(��Pc��G->���8ҥS;+-!���1}h}��Ö5�xM�B�U�!�d�z��CR$ښb�*�11�Ք�!��Ş��0���tc��@H� 4!�O;0J�� C�n�8ʇ��C!�䏂e�����m5&%k�&32!��S{JHB��D�M�����V�!�[�F���&թx�P�C�1!�$T�$'^��A�ň\� �s!��?$!�D��u5<�JG���qCp��cʤ8!��%hK&I.d�TI@�E g7!�dɰ@*��[�(����_�X(!�DΩ����@���J
(��gN�c�!��3딙�ѣY�2�"bf��6%4!�J�4�9H&�ۚ����F�J#U!��Rx����HM��h�!��5V!�Y�^;��;��g���k����!�K� dA��ėY�
�1��R|�!�ė�`�<u�נ�y��ђ��~�!��_���%��0�	J"�U�!���6��-�b�{��85A
�j�!�dU�G2��z�l��ǌ1	R �;w!�DE&~/��
3a��J�`�,εS!�$T3rƸc�Вx������#W�!�C�64h�L
 b\h`/Ư}�!�� `�ۡ�L16������Sl��6"O>HA�A24�)Xt�ڄ\�(�0"O�x��Z YT��6LL8�6X��"O�uS"P�F����]�bS\)�a"Od8k1�@�{f<YG#�\e�Y�e"Or��v�
3E�$d�P�,1dtX�"OD��LLצ��@F�C,�t�4"Oʈc	�� �-v�и6�lPcc"O0U[���j&y��c��J����"O�<�p�ݞJ/��bCaɑo��0�"O� #%�S�L�5��6>�X7"O�hq`+��,����D�^�j�"Od�3�((�:���3-��9D"O�I2a�6C�. ڤM��oN�{Q"O$5����:��Rvnb��8i�"Oƈ@v�ö.�� �)�MP�?D��0$#<3�.�y�JV�L���>D���p	�7pG�xq�Oe�DB��<D���#�Ѱh����w�[�VR�l��/D��5H�Bo -H���x��O+D��Э�=l���T��#`N���+D�jQ��)LQԨ	��]�D#'D�Ts�! �j�*���]��h��(D���'�'_{:�-��Ԭ*D�'D��0�	��	�ݘ���P$�t�E�#D���D��(�f�K��>#��t�=D��r��c#t�82h7ԀdCa!<D��
bM�8hdZr�ܚk�j083�-D� g
 �nC$�:d�Z�i�<ԓb�,D���5K�!	��4�ř� �rȶ�+D��ГŒ��L1+ ��.�n\1b�)D����x	{��"c��HcH%D�pbwǗ�w�2t��'���R�>D�����T���`�%�_s���D;D��*���-v���J� ?H �h��3D�hز�"d�
��r�
v�葂p�2D�$��-F(�*a
@��cN��5(;D��`��5}@8��
H6c~,�4�>D���h��V�^l+���s����H<D���
5"D�[�M�_ޙkvg$D�x�HC�P�=�DB�$=޲�j"D�#��<\ĳ��N*	5d�z�B?D��ꤩ�4"��u�MQo<=@�8D�d� M��8q��f8q1�G7D���e�6�(ف�J4w���"��6D����! �A��a2S���v�J� !D�|��(JX�H�À��\C2��!�>D�LH�:	5DQKr�O�7�D�#v�'D��k��ݕTN�aa
�	�(�9F@1D��`F϶� �� �f�Q�B-D�H�v-�_�<$�1�@�(�p͡D)D��S�P�/��y9�o��3��41);D��+�@�Z�ec���A�d�)��<D�����V��O\��2t�g&D���t�2��U:q,�$C�>劗`2D�H��XlC"͸�˝�-�9�a-D�����2�����_��У�J'D�\�a�*E��:2�*n� 5Hd#D�$�d
2 ����̡�J	�q� D�x���#u��c����$���"@�1D�� ���}/�	��ήIނ��$-%D�$1B�I0�� cK�AцЫ��(D���Ƨ=w�p�%�E�m����N'D���3�4'8��'�L��1�$D�� �H�j�K�Q��^�5�D��"O!��jِ�����
d���"O��as�L.&�T��b�0��"Op��B_	��e��C� |����"OJ�[T
��`����y�����"O��:�N��o}��z�"_�`�� "Ot�{r)�O���a��]�����"OPͣ�l��I��م�6�b�p"O��y��K$�߆m�Zi��"O�������0���@���0�"O5��t��!S�&������'�4`��&ԧI��
�`T+Nx�9��'�ک�V@M�'����H�x�z�'j�!���	������ݓV' ���'Ҭ�j����\�=zt酎K�R	;�'�\����	��ezc�	�>�4��'�(ԮF,I�L9#jV�:;R�j�'| �vk��4bB���3c��X�'-`0{ECu��@bh	.Wξ`:�':yZ���58��@�Y&��	�'���kC%L�[N>�k��R�{�n���'���kL�-��u�3h�1D��+	�'H"eR�Ѕ>�D��Rń�6��)��'�ލqe^�+F��H��T����'#���c�O�u��,�Pʔ=��U�
�'�>�B�n�f��IQ� <q�
�'�а @��
���
�Q����'�F�kŅR�5�~�y�	���b��'��(�Wg�?\�$�"ra�Ҡ���'�D����>'����k�a`0�'>2\���[�4a��A$DJ>{L[�'�}�pG�W0�����ե_sx%�'\�z�g�Z/L�04��"T3��r�'��
s�\�"!�	���8Qb��!	�'IVZD�tߊx( BΎO�>x��'RxA@���]���G�I�]��'jP������ĕ[�/IF�r�'�Гƅ-zJ`h��N+=�~P��'րP�F풋,����D�;_+X��'|�=Kg#�<�xTr)T�Ic�:�'����tM'lJ|� J�H�����'2x�*�V+�T��h>4r���'�&t�L
�	$R��5���;!�'v@)��(t|����N�8)h8�'���3`9��l.	�CXf�@�'/B�c��$I^���N�><�b�'�ʥ`� �0�vh�s)Z�0:t�A�'�L��%S�0H��2f)�.2�h��'����"Ɂ2uB����h�8.a�T��'��1���B*jӬH��"��"�d�(
�'�x����ҏ8Q�P['�»,��	r�'ː�R� ֙nJ	����$�#�'#`���0|�L���] UZ���'��,iu�F�S���')6���YD�<�b"���7*�A�^��bjWu�<Y�C�t����v��{����V�II�<q3Ʉ�-��șRK�u(Ő�,�C�<y�b�.V�i����H*�)
gJ}�<Y��N>eLԥ�s�Y�}�4�����@�<!��2@n�J��� kB����LR�<� B٠2!�y萏5��m�%*T���Q	]�k�,�5���`�h�aA9�1�O d�a@	pX�Mk�@�]�ҕ���'C �n
;�Vܙw唴 �|y��?(fB�)� �Q���ѵ�>�����p���4�'ﮭ����P�����A���;��8|(}��Y��4)Dn�sѶ�ˤ/�,lb�M�ȓ �q��G�ݱ��R�.����ȓC��a7iI,�vD����B�I<�H��	�Th�@��[�zֺ�����B�<�#ǟh�R�9���k3�B䉿>�EbU!�S�8���@1;����$�"���f=�e�K�%M���16`��p��bH���*�'����fnN2+���=�����$�P?h�@��/�R�j����yB+O�
&���&(��qA�斛�y�G���{�!�*K��IP��V0�y�g�H~�!�JQ�e�a`�$�y"N��2�Pz#�_�R`��.���'�ў��,uآ
�w�d�S�]*3�
�"O��hRQ���2��Y4~zXr��?}�)��3�����O;%p9Q�@��C� v�$2`F���X�kv�߿y��І�I_��R��L�A�P�Ag.������d'�D��xUI�M���2�Ĕ4fQ<�5�9D�x�$�����r5��B�ޕXB�I�vь�.�����	��[�j�pB�	'<�R�3���7{�5��K�~V�܇�I�HIt���iUer����G�-r�>B䉱e�A�!c��B`�[�܇$<B� kn�ءo�<AT)�'G�Zo@B��If��E�r��-ѬP8"<ϓ�:e���+��T0���e�VՇ�@k�iZcb�4Y���U�E?:�rm�ְ?�2IF�zHZ%����t�N�c���<�N|j!ҟ4Xq�g/E eJ�)�c�N�<�2h��/��������,�S+c�<aU���	��y�+^�h�x��\�<!���[FL���ɧ?���8&�U���7�Ӻk!
�Z
:�H7�9�\B�d�R�<����U��m��L�?\�ʂ��P�<�4B�.>j<� m�9|�y�P�<Y�K��2�m�tƜQtf�Mh<Y�� 7L\�y5&Z�ˌ��eG �y�(�>BR�p2L��̤²����<A�d��[MlI�V�"0E�){E!�$9߾-�S��)f�*p�Dlc�'pf�Dy�dƹ��	'o2��Q�`�� �,��ùc?�B�	,+&y��
¿;��bf�\"<qa�	]y2�D6X6z�ш�	C!ۤ	V6�y2̖�l2V�R(�$��t���y��]`�p�ku��<֢Da�Q��y�*F!vj=#�gL,>xUbG��7�Ov�=�O\�@�W�G�)����kK�fi���'/��aT�D�4��8c�_[� 
�'��H%���Bbʀ�BuT�c�O�=E�b	�h�6�悈 nv�3eJ:�~b�'3�dy�*P��Ճ�m�0�\)�J<q�
��I�	�x���۸�Z s"$�zE��$*���e�W�1��r/��4��`�f %�a��#~�%� �Jrl�d'˲bs���OP�<Y&�#LV��+Uɺ`A��\I�'�ў�oq���("��� p�Y-'��ԇ�^иS�`ߩ����ħ̡��l����a5�ݫ%�F	�7gY��0�ȓ7ly�2g֒T��E�0AZD�b���_�MR|B���6zl�#�M�d ���Fd���@�ұ 8,��H�-��>Q����� ���DmO�@�T0�MGt�PY�"Oj�14#>�ARP�e�4���>	)O�R��Y��Jvl�m�D���
H#H�(Q�C�?D�Ij^*"1�T0ISP��DC�}��C�	.4B�y�̎�{���۔@�>k��C䉔[Ŏ��� J��fAK�'(����>��ʏ�a�Jaq�LM�/��l�t�V@���'��	�<1��Q���cXZ7|���D~�<���6hʴ9uO���U��(�v��?�J|��&�6yl9���!"�-j2��z�<����%�8�R����j��P��i�R�<�B(F:�X�ŤƑ�M�O�<�!@��<�Y�b�)jJ(�Ј�N~��'� �y�O;,ڔa�cd~�@	���d�o�Zd*���M����ǳ(�!�$�~���#�ʰ����ߙo?!��:v�L�Z� ��$tę
c�U[��.�Ot0BbN!�N#!��?���I��iў"~nZ�thE��b9p-��i�+0"?)��鞓F���)�+�
iu� �ԡ�D3�O��B(�`�2�1�&�F����"O�!�(�
B�H�f�3rJ� �!�D]�B��X�1	D4�>���!
�2�1O��	�����'���HP�&J:T�f�0@��%�0?9-Oy��H��"6�e���-Q9��9$�iUd����dퟱO��$�B�������=��-��D!�䋄/>2)i�
X2z���J�l]!򄎱-P����A�#}�A�P��!\a}r�AyB)�F���6)��}������hO����$�]�P�
q�����W��4e�D1�S�S8>�&0tނ\hp��2`\)�*c���I?TN��2 3�eQ��<�7�͉��I���x�%�$�p��'Sr��Vn���p=��}"�S;I�Q; GŒR&�i�f��-�y�P�Z���M��E�R�:wA8�y���	��HD�T�r�D�F�N-�yB�]̠��գ�p�2���-��y�JϠ?Z�P3PO��a�X�1����y2Á%	�!�5��<E1D1��/͊�y��X�2��MCv�&��衎W�y�Ì�fA~�cEX�PJ|�!��y�!'
M�0̔�{��4x1j.�yB��8W<&���'��<[����^�y�����T*e	�~9��P����yRM�yd5��(�7z�!hw����y��O�_��X��[�����v�Ѓ�yB�#�J����̥�T@���y��<t���يj,�c �7�y�\%���B��,ꑏO��y��Y���Y�`����Va��ʡ�yb	Jf�8�f�h�ʴ`�]�y�'͟-�H�����*������y�'�5K�=���X��F$	�y҈P�lS�x�$HT�]i,@�5j�y�',0^�%�i��S��e��8�y���w���� yz~��1����yR��'I]�TkփX�k�5[��=�y��	O�(�p`�;]���#��C��y�
{���3��O�T��2�
�y��o�����҇^9�ȱ��y��F=<]	0��3P��5[�1�y�
�-�ʁ���H�}t�B�	�y��6{7��U&���p�lT��y� ��e|���`�=��$�����y
� (��dE�9�>Qc�2g��� �"Oʄ�s�O9�ʐQ�!Q�u�zu�r"O�(xlۺ&I\�U�0ٔ��"O8��c��VҰAkр��&�4��"O��#�B�L�i�O,}�4��"O������yhZr�MI�V�&"O���1���a$�r1���t"Ol��C�<����fe�=���@�"O&8�T�T�7Е��M q�h ��"O��RB<J����S�B�v�00�"O�в蕟o��$���Rüi:W"O$���O-?i�1 
�&�,X�F"OJՋG�I�r�|� M�IL���"O���U���j�­Q�M	�iB�5C�'����a�,�����T9,,j�)�C:���'��Ps��{��D�!$4��X
�'�PK�n�{�R0H���	�@��
�'��cF!�W�6$y�eܞ	x���'X��`0h�,H�H -�rnf�`�'�&,SV��?e�"�*�ޙsa��'9��xAŇ�2� ���qU�Q��'��1�3
47��SH�(:q� P�'0������]��(�")�?�p50�'�ݻ�o[�Lc����ʢ(?���'�n���+%!����m��vfj�a�'�֤�E�?
ʠ�I
QvU�l�'���!�b]��B����/n�F�a�'�������m��]ڲʉe�d��'4�eۆ�Z,yF��reħw��s�'�R�k�	ىAð�@"�ڲ�`���'攉�@�j���G�� z�'(ɩe̟�Q#�Ջ�'�y�z�s	�'�ăS��&v����+�èx*�'�֡�B#lӦ�1���"�J�'�0�zQi\�^�@is�v�6���'P�PIP$�Q���Ctϖ:���H�'!�E�r%W��n��#�x��4��'�Ӗ`�
O�d�kR��)D�dUH�'\T9�0�G�t�z(0Q��'6`�q�'��14A�1�|��,��8<*�'��mk`�S�p>=��l >�P��'#rI�'GK�V��C3ꀗYz�	�'x��P�Hq\�9rĞ�Xz��
�'&Vy��8re\�F�L ]��R	�'��M U�4,���`�GB�J\���'�2�3lޭd4�"����Ɠ�y́�j�yfu�t���yR!0{1Ԝ�F�[�D�DÞs
�'��<��h��a\"|�� [�yr
�'��C��_�ʰ�A��}c�L�	�'nFE�3C��C4Bm6�W�u�^�H�'˸j���8Z�h�F):����'oXR6�J�_�
�ɤ�N&8{�'X�d[�Տ6X��JF;F����'l�!�+N�Z�܉0�[`,�C�'8�􏎀�0(��W
�b9��'�~!���	����d�V�!���	�'?�h�"�7=�a�S�֭T5�I��'D�ШR�z<�A�''Y�C��x;�'�5���%�)�
��J�X̐�':̔���Б#��P���t��ѫ�'�������0��!�P�Zd�u��'�D!V�*w����7D����'�l��Dʖ])ԅa��Ҡ	�&��	��� z�ǉe	*] !X�p��S�"O�q�d�5޸Epb�9-��a�"O!��KD�FT^e� ��W��\@3"O0X�6L�'H�x����.�x�"O��ju��=c���{�q�J�P�"O��
!	�r��@5	˫ΆɀU"Oʝ1f��9���jL?I����"O��Q�	�>���w.΍��4�"O�u�`����.�a��� �<�`a"O�L8���%l:m3 (��
d(�ї"O.=����,S8�(�j^�mXD�0"Od���r�I{��1; �Q"O&��E�Y�,��=�ǧ�)i}4�{�"O~��k�<󰸣R�FZ<�R�"O�|�ϸ6��������9�1"O6�� �^�U��(��H�V��""O8��Qe�����"B�J��%�"O~,�E`ξ�@hv�Ġ�|�I7"O��qF��
a���2���C�`\;U"O6���NШx`�����Zd���"Oj(��O�U�f8L�.I!�P�<ɇ��6����%m-y��1g�z�<��ɔ,b�̻�ņT�t#�v����9��{�� �7*����EC�d�!!��y��4X�%r��
�*���Xf�֨-i�'���p6֩��Ϙ'�|��Ĕ99��bKN�Ai	�,/<�c&�Ŭ����Eڣ����3?�ܸ8�(�[\�52	��l��y�!��g�x�	�BtGx��l�8 ɳC>X�"�pe2�
.4~tt����L���N�I~!��1w�*%�
�`q��]�Jg�C�I���ʽ0ь�U}֍�d�i�q���9�4k��(�0 �.��dB���g�V�<q$�����[=7oP�Iu�J�6��t�`bQ� &��C��U�R��(A���"�%�,Q�;S\��G���� �'��a��3�1����ZUR9�a(�p�*�N�/j�M9g��_�8�'`�(���J�t`s� }��蓶M��eǘ�ҦkJ�n8Q�H0�ɂ#-9��-Z/o���MV�<߉O�!Bg�9[��D:�R�,RT�'!��"�fS4�bm��I&n�BN�B�`p���4 Tp��"��LJ��%jo��I�)�5r�0 1iۣQXz����R"Q�p�� E6^�P �' ��;d��= �nѱ���?Z�)�i����$V/>nl���
> )�_}H�y��P�K���YD&��
06���N����D��iV��Po��M�����W�!�AٵnUB�İU#��S�t�:Ђ�^�R�'���F��{�!���OLH&�02_�FxR��=A��s�j�7,�����D	gf,�aįrt�qA���~B�ޑ)j�3��K��XHU�r�d�DY(?�>�Y`�ͥ0�RY1�떟HC����c��O��(��8B��dFЪ2���c���<=zuE� u��=�ȓ��H�
L�S�Τ[�凾B͜Ml��V��7�٘v����GHٲ��%��(�X?y�Eǿ@Ϟ�0z眭 %f8O-�%���/L����`�h�C�k�����k��W4/��M� @�
���H�G�.zp]��|� �O����+E�߸��	Cg� ��L~@��U��Zt��2��.��Æ@�	vd�}B�Ɠ�l�
Y[�C\0P\nhA%C� h0���&:���Ē�,k(�蔣�Z���Cf��k�&��2�C�J14q��J	�0d�1�_>���ŗ�"�Ԍ��X�lg��l��M�Wgɽ=ۈ �f�<D��)��Q�q�2��F �-�d�A�S�}"�BhV��i",�!M����ҍC2L���5�:M���_(�"��Q I "����ߨ�.���`��'��Mcj��j�#�Juy���ƚoJ�]k�8���7؀���Bm�3}"�
�0���SG��r0,p@��r3$d;�%��h��PSS�:v�  O~SD�C���ȓMؐdłD9�M��IAHPjĎ��?݀��d��B�5�G I���ɳLQTq���$ې^}�(�$*�=�eieW>�S���%}�<[�U��5il�6�q��(�,�Մ34�h2��W�H�����LB%�t�X��vI�4�N��8d2AAȧ1��#I>9a��&3��ϧ#��m�U$��. �"PAT�D���/�b�g@�R�^$c2JiC8u�-T�	�mI�A��<�V�3�	,ND����IF�	s���"sK�@���B�j�*\iL��P�	�G��q��W"d,�z$	�?Y8t��żCF;q�X�J��b���8V��OH<��� �:b�ꀈ*DϿMʼ�D�%y.4�.�*!G��ˤ��N�2����i9?)��� ź�y����lqp5��d8��F&A����Ŝ�P��HD�r�֥��B�&y�-���K�N|�3f��g��Q�@~8��rB%M�(�Vq"I�tz�`#�.}b�����(C�ƞ]~��� &��A���>>��Di�Ծ��XC�Å0��=�`,�=�L�;�RY�ƌA3
�Q���M L�ÍE��I>�6(���+ޒ!H���O��C ���yG�SX�=�b�� �<�֍İ�Px�	ͭ���qF�X]�8$LC�Mς�Z��=e4 ��E��B��lH�����CA�Y����͐n���n������7Ob�y��K�i�Of}�vgJ5EL� �o�tU�wlV7kq�|��ŏ	���n7<Ol�B��&6`�ax��L�Q4�>Ѱ� 82�0�( �DAvh q0� ZF�P(��L9�����}{n=�b�_C�<�S΂5��,�"�,Xt���dF�= �(�O�l�q�gwD�I�����B�S����B�@��LӰAπ
�E*��� d�!�P����`w�X�e&�kf.ψ �Ј���q��ݤO9��c���J'>�y��P���pw2����<ۺ$��qu6�	Óx�&U�Gr�b�oSYhj�x�ʓ6YiV���d�(�:U��n�]9r��[�,����ɖ pن�	:
�&9P�� ]�$�iW��	vq�p*�MA�"9m��$��d\l��ē@P�XT*$Z�}C���")�>i��GJO
I) �(Zu�`���D�8<S�Y�#^�l|Ȭ�b��y�ɔ�n� �+A.��f�" vE��FÆ��?��ER6���Mc��>�6�DS�L3.ڹ�3��ib�C�#zۖe�SaP�2��T��ə�@9���٧>9c�L~���9d�9Ol$�4%�
����k�$D�1A��'����I��fF���Q`ӗ+/>Lc�ɹ�z-�2��!dpH�BCt<�u�8n�RC2Ԯ'B,�U�FkyRLIQ�>� ��V
�nm�T�*SȄ�(��)�,���dJ�)�B�8ą�,V%!��߾%�`,{$H��Y��KD"F���#��ǱB�ġ��{�N0J$�����)�z�d���S�E�?�b�3sN�nO������/����7OD5y�P����&��`�ӧ5�J(`��	�6]����%c ez3�'�,�A���^(b�#c�H^�ys���R'T��%bW:1��AE�5t�"�yD���E#1��!);6�Z0,��hF~��	�'c��(��a	S���=D�p���'#^iXSș�{�=��+O72�^�HD��2���>�ʵʐ�o.8�G#0�ԽY��$D��
`�+4y6��ԩ\'lhb�$E-b�j�'9M��U�v��"wC\�O�0��D�xBb�?9X`�a��
i���F+ބ�p?�g���/� �qb^�~�d�D�WO'Z�0�AX1+����gɖJ�x���0Ӫ��Ҍ]��VfِQ.Q�t!S��)��=+��NP�M���jU�8Eh����Ok B�ɶ+"��#$��h��8��4��I!P��Y�� �����h��R4�W�vL��s�R�VB�L�r"ONe�ȏ�G���B��U3���re�4}�ƅ*d��٥�(��DQ��nt����K��=�/řuh��Ѽ	�`�i��Y>(�|�q�; ̈�BC�'+!�D��^���TDA���M���%�!�_4te���Ό*�J�r%��>T�!�dӚd�"���Ɏ�g/
�I�H�!�Ĝ�/2���)��Qm�i��7Qv!�D�M��uД�ϩ;Q���VbA�ac!��Ȟ|�6��.3+j�Q⊷Y!�$>� ��sg�>s��� ��!Z!�dF&�:I�����[����ѲHH!�B�O����w�_�]��HX-O�!�!�G4$Z��&g��Vt랠#!�D.@<P��a 0hxl�fK�(f!�$��,��2�PMZ,����['S!�D�-�� JRh�sD��h�^�(N!��!	*���	��-�dj�5:!�$A=w�TA�cq,a�N�V!��S�.�pQ���=fP�S�&H�!�d]�L[~��)�0g4,s��޲&�!�D	�g�6�6.ځ7�9hע��"�!�$݇=�88� �
2z� �bʄLc!�� d��GV�����ɸ|~��"O��bÇ����.ګK4��"OڕЅ�H-
���l��}�""OB�� M���{b��
Q��TX�"O�݉S?Ԩ����E�WM2�"O���%~p��X�/X�T���c"Oz�*](�����e;AKǮ[7!��G�A���D<�yU�(Y:!�D�[�$Z�+ь��F��g�!�D"\�{f,�+3��=>�!�D.������٘�|5W�3[�!�D\7$�M�@KV%3�X�$��k]!�$)J�� 
�K�}���{��ٙvo!�d������K��9(�#q�̀SJ!�D�-Y>���<DQB�ǐ�+8!�T�:�b gE�g�!s'皪G!�$�(.��Hҥ؛���af�;/!�
91Kv����3=2b�`��<=r!�d��g����|!|y؂�X�!�D�2&��1��0L���*$e�!���wl岔�^����:�!򄞊%��S�I�<�����!�ęK�*�z�'[��|�ŉ��I�!��J�Bj���BS�+S�a3K=L�!򤁢@Z�X�U�Z�KY�h{�$�f<!�DGx���E��Z>a���^2$!�D�7)z$ВB��^C���c�!!�dH.{m~=bi��9X1ah�t�!��ۻuQHcE%��<
�urm^�Q�!򤜾BY�5BB��+aJ����E�!�dE3�F%�æY�p��c�P�9�!�D�kQ^�srgQ�X�,�)��D�!�A�F�ӈ�6�Kx�C�I3nx��Jp�h����T��$�xC�� D/Dݳ�!VOͦ�9��_10E�C�I:Rb6�2�:��4��ڏ8<B䉅,��=�S��/ǌX�6�G�#��C�ɿx�T�2�� H����*j�C�ɪD
n@&�KJ�5{5OD�gs�C�ɐ�	3dƘP�(�P��)y4�C�I�kԩ8���c�����э-�C��r!+�K�lʤ����R�F}\C��	o���P��O�~�b�Є��{w�B�I�wRlu����=\
$ ��G2"�XC�I�,�6ap�d,�>�ഥ��? C��=, $쪤��I�"h�G^>M{�B�I�B�(��?[*���-PB�I u	(�k����F^�=��j�^{�B�I-�	�KW�Dxj�K�׸h� B�I�e��ܠ�H]V�N�	A� ,i>B�	�!r�t����bp^�S%F
�6�TC�ɞ;V�9� �5jbi*g��f��B�	�i�b,��Yz�x�K�;@�dB�ɻ\�H,ۂ�R�*��c�� �bB�	$ג`��BR���raO5��B䉯�*Mb�-�ri�Y�A��$>�C�ɫv>�5 G�V�6��-�`��~IdC�I(Y{T� Њu��o�2�xC�ɟJ��� �VA`5�Ҡ�0\bC�ɞ.��m�w��.���)E�X`�@C�I�c����tmV6x���#v�@C�	��R���'^ �q��a�hC�ɩ-$
=��͵s��B�$o�JC�	A�u��C�5n Kf3-aNC�)� �\�v��	Vv�0G"O5^^�#"O���C*IuAU��"_ ٣�"ONq�C"�`���y��	����"O�`	ՋۖN����e�m��m��"O���ÇS�����MdLh��"Of!�%įt� ��A�� d9�'Ĝ\@��
6⸳�MJn��Y�'��(xWeΦP6�x���[��*�'��X��G�i\Ĕ+����o�f0��'9���֋��b�٢�ԩe���'!p̩@K
�K$>�*���v�
���'�� 2�εU�v�'�y�0��'���"`G�[�(���qs��	�'��љ�m�=�F��v�m>����'�l�WoQ+h�t�H�臔c�`��'ڴh��G�g.X{e�������'�\�W�O;`�P���9{R�s�'ƌ��j�,��t��I�h����'�Uh�F��Z�&�z#b�!kQ(���'�M{� �� �>y+%B�5����
�'�\P�3��4>��2�.�4;�^��'v�I�3��
xlR�Ka���� �'��Y"��3r)0i���ru��'�� ��Ѷ\�Nu�˟�q���'�,\�uοK���� 
 ��Q��'¸k3a�kVz�J!�F� A4{�'�|��� �8#p�M���SM�t:f�B=*�qO��� ��?
��!M'�$��"O�`P�k'a�&� 6s �� �1�� 4v
�� ��7K�, �q��e�V9�cO���|�d=@<Ps��>c\�� fÿ{�
�:�O��PdjAEcaR�r)����S���Q��GB$HDx���  ���7u%�8�$��4_��i�R���Z�쁭�!��S�d�"ȉn��o$X��*+L:�{V�B�;�,�7ƃ{��������T�t��4V[쬳��� Aj�۵D�%��ȓ��]qsd��� =���$n����QJ[5A6�i
Q�jG�}�f����Aq3D3�Ď��U���ΤT����Fݦx��Qi�(�i��d�׉�P������ϧ�0`�P�2`�z��̑[��Y�
�� r<3f�a����/N�?�d�@U�L�t 
"`<�o\.&f��ᵄ6Iѓ�S-�p����df��N@ĳ��P�)8�4hA�1�~"�<��e��'�K��,b`��9
j|��n�=�Bp+!���,4�� &G3?�^�ۑ��7��>��f�Z
O�-Ai������V}���K��"9�!�$�*��-��Ȅ�M�}���B	�06M����1I�I� p�"�SlAS��0}b�����Z��$�:���'
��{eϗ\��d���9T�p�	&��z��E�$�"���0D~P�I��G�--Hd��o�D�(�REՐrf�m 6NMB��(ذaӝ�O4d��ʫ#��t��l��1���ᡏ��U�ࠫT������O���Gܧwǲ��~��L�v+��+!ސ���?�<�ǪN�m��<�b�(k����S���)i���� � }��H�`DI�blrgϯ�\�(�-�|�<�G��h�t�kgN�4�Ƞ#FE�ɶm 9�Q���b�+T��n?a#H�8`����h��O�S|��L�?/����M��I�bD$:r��e\�x0�J��^)i �"�~�b��
Q�X�}�OZ�#�/�3.��A	S��%d��I��O��1g�'Y��	�g���JivB�0ybU�U�ߑ��>�L�\4� ��.Ϣz���j�)<O�4�w�Ρ|���z�O���"�	F�����x0f��0"O �J��K+&�������Z4jB%�|�X
_8t U�j�O���+0'|�y;��$����'��	��V�x��N(�5��c�j�'Z2���>�s+U�x�����T�+g��21e�Yh<yЅ��_[�R� �GzP(vMȣ"Y��\"D���Q�i� =�'�G�'ֺ��TjοY9�y2��$Ѵ��*�}��	=.��Z��aG�\P�%�y���[K�[ CU>Q�x5S��Z���'�|%{�Z���?� 4m�DQ��8i��*6V� 9�"O�b��E�U�Ԉ�ĩ��JtVY���(�qO.���Y��;e�(���Q��
<zƴ��:�'b^�P��>�%OR����ꑔo��M�ACuH<��+�ɀe+W]T8R��P�R�Ƭ�n��p?aU���Q�鳆��*`���.�Q8��*�ڇA���BЛ�DB�G��?�4q�,TB.��'D��B�@>p��}z��՝+�6�g�/}ҀK�?]LE�wN�_�:U\e�^?Y���G�5�����+V�IR�&D�x�w��" ��+�"�EiX[tL%{��'�ڤx&��M���Y���2�y��V�%�b�����JTp�0���Pxb9�����ōA�2����G<rTr,�Kv�RФO��p��V�5�����d�/p޵���A	x����<	�x�&�* �5�[~~b.�>V��MQC�t���vFט���SEHX0l4�Q�ÜL�4�J>Ҙ��A;L*�Q�Ox�SiN�s�X0�L<a�R��$�h�'�$ �bGx��8#Ӯ	n\ZA"�'B�Y{�lL�.|�`�N2}D-�C�5���g�.�bI�i��8��u(�Do�����R����*1!ҥ"`($��b�$�>l�h�)樅�f���F�̋F.֟��I+'1����͝-��gy��G�pl�Jh��\lY��e�0��<A'(�]nO��z��M�KN�B�j��r�Z��ԫ\�%>������-�a|rc�lT��M�H��@@��p=�e��n>x'U�v0��t �F�p�a�G�#��A�吊͐x2	�Y�TP�Э��}��lF"��'ޠ1����%Vb]{�C	A�q��uB�FW/��E遯��b�>���"O�ht� ��oH�4��F�	�zĐ�α/���[#�i��#}�'��=�&@Z1Tg�A)`I�;1���"�'�f�!�ׯ�P�1� �0� t�N�v�Bq�p�[S�B�0<aD������;A���⃈>o�x���N#��p��]��� s�
��*�� X��T�&g֗L͢���'�Ш a�G[�8��Y=XXjP+OeQ���0f�nIɁ�92 N0�VGP�7K�c>�j��-�tK����q��+D��w��t���!E�N��J*F�x$=)�Șt]���I/V�l�� �o�R~�%ԇ_�3s�74�5+�gĜ�p?Gg��`�M�Z� � ElY�p�V�LF bԨ��MAVȎ�[�oă;�t��'4�B�J�Hz���՛[������D w����g�	ouD��5��I2�z��ضV�`s��L I����-ʭ8��ec�'I����";L���-�:���'�刡��;K$t��I�'����0�ю$b�>IaB�X�A~�tUc�]K|�`�e-D��*��3k<VHP�AQ]6��%�-0�T-��#E��x%��*'T��O��-X�x���<�L����Cn��s���p?q�T�e�T�Є���$�)��#7v��	�IK�V,9aB2J9����D�4>� ��U�͉eE�;:Q�|h �BWx�u�^\�S7�ԭ���҉�xd��K�dI�B�I'G*!J"BѼq�$Z���l��	�ꑫV�;g�$��h��41P�ߔ!0�Ͱ�+��:؎ȉ�"O��s%�Y�j��j�3�t�I *;}.�5e,���@4��$	�'�t�)���C�>Y!V��/8��n��&�xq�͔0"��\��)��<�P�̗7,�!�D�	t0n� ��{�H��g��M!��1H�I�EX�Aް� ��"F5!�˚>�`عCJAIa��D�-8!�D	�J�����2CJj�́. ?!�D��F9��)w��T؈��$.��/I!�$"xn�Ix�*g��g��OO!�˜L�P�Y���*����f�J5!�$��?VL���mDL�����eE�!�$��b�J��wEGsL����E�!�D�C��Li��9�(�S� ��+�!�dV�$�<��rA6#Έ�󥏠K+!�d�5W����o��D�v��ꊣZ!��l�F�0�U�o��e9�ˉ6�!�$\-�(!6��4B��%�#ʝ]!���v �4k�)��y�.�Zu+��.1!�� 4��e��H���z�
��֥H4"Ob�p!OR3Pj�02�ʉ�[�8S�"O��� ��r<�4(�,�*���"O���G�!h �S��`Ԯ486"O��y�bX�$S��J�Jϡk�Դ��"O�S�35�(J���!�����"O`!r���{�����%�	-yTɩ�"OJI��D|鲢��wv̼��"O�̙�`��?�P͹�		cp
�e"OfA	��ܛe�r�Ȑ��p��y$"OT��!k����H�+	?"�Е"O�)�燔$%���+$��xC"O� �'��l�-:ԋ.�"x��"O�U�B�<7��J�1��@҅"O�UP��T.�0��6&��ԁ�"Ob��dߗC�ͳ�/�F?8�zd"Ov�����Hб�nLp�0�"O�d�-`Nԝp����x�@�}�<����-k��Z�D ���r�
P�<1Uh\�A��DʷFK�M�i②�w�<��g�B���!�	@����t�Qm�<y�BP=D�����?V<a�Kw���#E�x
���=/�E[u��3U�xt���2D�D@b�O�~�vi����Tm`�'1D�cgH�|@z��!��3DR0�)D�$qs  �x�0��ͼ8{f��$D� j�b�< *2�9g� ;�,� �4D��9�L�	"8�Iw� ���F1\O� ��ԇ��,�d�`���bS@���A	'϶⟢}*��1I�N����I�V�]�e�2\� ����IJx�	ېn8\	�g x�2�סC!����C�@{С���M}��t��DC�g Ȁ�Wi�FfX3p �r�8ZF���d@(��0��V� BY�nY��b �'- �3�ɳ+�� ��:�j���hſA��(�,�S�b�$3Y]���h�0|���V�AK���OY)f�����<9��_.���B��n~����}a�u"@�*23b��rH"����WF\& X�s������|��I�g0��ԁ˓a�:i"�!H9�LH`1����L�"}a��F�.z+�t��!>M���4�bol��O��ۅ��$ �֒O1�ne��˜VAȽ�ր�%���{���[�48���nM�Y]��'UQ�4\>�e��^��3�Ę]���bJG Y������3GB6��0WD��Oq��7�)T�X���Y��'*� ���Q�lJ���Mߝ�M�e�?�j)�ӭ�|�7��-4�x����<`,@qjD"N80�b�
׸i�3���N4���O���Ո[?}�H%���١Jy�ش|�a���F�^!) M��O��>�enN�U� s�@��^�%��(��y��՗S��	����!'`b0�CC��y�#Hs�1����#r���y�b�x��庐eJ?5&��B��y�d��h p  ��   �  4  x  0  e)  �4  �?  K  QV  ma  �l  [x  0�  ��  ��  ��  ��  �  G�  ��  ��  �  \�  ��  S�  ��  d�  ��  b�  ��  � > � � � �" 7) 3 5< �B L �T �Y  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9��CZ���1.*��5���#D�������=9js����]>+-B�I�L,����ơT� *S"0G��B�I�<w<̉@���R��Xrȕ(Uv�B�	�n�t�hՈ7Cn���ӳ;�B�	x�Ψ3�E�V�B�ʑ�ޕ-bB�	�K��� L0B��h�'��O�`B�I~����b��L�5��£~�B�	�0�dq�  -Nz����� 9�0C�0>a1%
�y�N���.M7@B剖+($�w������Ο&|`!򤂰V�dS�D�
��PZv�I!��"���㰁L5=�����	�!�ӄA��a Q�&�ʀp`�0#&!�$\(�����N*�Z1�f��+%!�D�J�ݨ�H�UwP5hd�	!�$C0�d��#��1a��ɷ*���!�$J�gÔ�[��,;�2	:D��J�!�d�c�\���HOOj��q��o�!�R 5rZ@
T�� ]VH�RbY��!�dI�{g)#��MF�EQ�J�7_%!��= G4i�� �<+������5�!�D
�[�T��"D�*��Mr�N�2w!�$�aFڈ�&�ذM�t�D��l�!��.a��To��6�F|��,	�v�!�DQk�m�D"��W���wN@h�!�X��1R�/߽`v�S!/Ìk!���/uӦ&�(__�Ո!�ǖE1tܙ�I�X�Ļ��̓�!�ԉT���k�E[*E������6#�!�d�zr��h!ꖰg;l\��cT�t!���k~�X oF>@����c�#�!�8H�Lk��7�Fxk��R/�!��Z�^l2��^ a���Rf�L�,�!�$�� .!���"S$�*�.��2�!��0BYڨp� �:8P���KȝW�!�*@�X�Oފ?g��ॠ_�)�!�$�P��+D����z�� E�!��  �!�O�M ��#Y��"�8#"O<��"��5Jf<a�AmJ-�Xt	U"O0�8��+��k�삓���"O����HM6��JB1[��ЫD"O \�!�Ðq����g)B�6 ,AJ2�\x� PB�P*Ybk8t H�$D�� ���'-B�ր]�h�����.8D�t;���w��y���qa����+D�����$�!��J�q�Ġ��k+D�D3U��
u���9��U����y��;^t�X�WJ['�z�22�ۮ�y�o�+q!���d�$H"��y�I�n}['zR������y�A�?��pDkc8d����B3�yb�
�x�*�Y&�%��1��O:�y��\�`�x�b N�����+��yb��,h��i�JF��aVl���y�eɊ�lcP%M�:mtU0�E̾�yb�A�U�͑�&ǘDc�!iv��	�y�n²vl6�!�5�>PVaC��yEF� U����Q0CB]Z2�\�yr��`�й�Z/���-�\B�ɸ$�q+�����X��BDz�fB�Ix$!Ra�Л:q�Hx�D�-L�fC�Im�^@�a�D:p��ș3&"Z6PC�~�"�:'HIպ��1��0� C�	VQ�!�)ǝC��3���G�C�0e�y:p"B* P��D�*͸C䉶X�J	K�*�$v���	�k�'��C�I0�ȉ�c��*�"U	�h�
�'�} �A�5ΒA��V�-�1@�'>|��"�F1%
��	�-4����'�^Mir"�#*Wr�Ф��; ���' 諁nÄ�̂e���k�'�j@{�a�i����b��p�����'u꡺�i�K�IAa�D67���'�`5+`�P�{��c���B�F��	�'��E�ũ_#J���ȓ΂g�Q 
�')�	�2�؉kQ �E�q�pU�	�'@l��A���b�t.D�s	�' � ���ʹu���:�f��o�NYA�'�@Ц'�u�����M#_�����';j��s��z:�yZ���V:j��'jQ`u��(&�%; EKI���!�'�:��i��m&�� �Ci��B�'�Eڦi���
PӇG�7P:$!�'�<DaS#��x�E�K-Q�P};
�'��0#B[i��S��5����	�'��p5�Ëi�&���$�8oD�	�'�r8�,	G%��3�6��h	�'xڸ�@�Ir��+��U�<��`�'�����8M���k�(�3�\�	�'F��c
ցn��9ܹ!G�	
�'�F(�A`�Nn��NQfS	�'6,-�ѩ
),�p<`1a
.&�H��'�=��"��'�,a�탸(�L0�'j��1._("�ݺ�E����!�'��� �o��yp���F���'�nD��K5�
iʶB&-��}��'�`Y*��C!;�Ⅹ&
�nlx�'�,T�� |>�-JS�V��bu��'0�)m�\��}��a�/P����'����j�uM.�ׇE�<Y�5P�'�~��JI�Lx���;¨���� ��x�@�� � #� $h��'"O��B ��D�2�$I�r
�{�"O(�$E��jX��豉�4_���;�"O�zW#��3AB�a�H�o�����"O��#�i� oD2-S��:k�����'2�' ��'��'H��'��'�9)�Z�����F�
�+b\8�0�'!�'or�'�B�'�"�'h��'/6%0	�	d;��3�J�:���E�'�b�'H��'���'R�'���'�X�G(�g��!sc�Q=C�ybV�'���'mb�'���'��'I��'�ʑ9W.�����0d ����p��'�"�'}��'���'��'���'��Ԡ�.�Pق��2-K�Y���0F�'�B�'"�'�"�'���'���'������щB<�գ��-��*v�'���'�'`r�'t��'���'���´Ҿa�>P�pc�`�E�E�'�2�',��'s�'��'���'�`m���:����G�p�8�3�'Ur�'*��'d�'\r�'���'[�YEF�!G��٨��$d�$8�W�'{B�'��'���'���'���'u��a��_3Y�b��֣�1?�u�����I���I蟌��̟������۟��dCܮO*̽x�A1	�N��Bϔǟ���̟x�	�d�I��������	ş�Z��澱�$M�x,̰�r��ڟ��I��H�Iڟ��IʟH���Mc�Ӽs�O�����̉�M��eLL�a����������Ц�á ��{1�8si;����Jl���'�b6M4�	?��D�O0qk@c�+jXi�� >FqӤ�O���Z9��7*?Q�OU��) �z/b��CgAvqʐ����)��'p�V��D����%Ea��c�D܂ ʱ�CyL듣�d�Of�?�����;��y��b�����VlI��?1���y"^�b>M����͓��9`w�\3�dq$�_RY��y�l�O�y���4�t����W:0���V9 �(� G��<K>�B���O� @�/� @@М�&n�-[ϜA��,�	���$�OP��d�L�'����\�N���h=Z/��8�O0�dg�v���iP��?�*�O�y*�íP�v0p�A5���PI�<�)O���s�<r�I�TN�2�*��$}lY�Dg����ثOVʓVB�6�4��|���,.����J�"T���70OX���ON���=|q�6�'?Y�Oy���J�aj����{c������.;:�N>�(O1�1O~�
a�9P!�L3:�ި�t��8�O���?1����]:%K�-�Q,�^��\ѧ
�&��R؛-k��H%�b>9f�@�2���/��X}p��KL*��|y�E@�z�(�ɮs��'���.���C�Ȗ�W7y��Ǹg=�����M}R�'6�БR�v�R bUNG�!��傝'�"7�9�I!����ΦY
�4
��j�3�D`�#سy�<x@�Lr�� �i��O"�R������<���ֿc�̉'i��h�a��-W�V��W���<��,�<�� /&aڰ2È�����*O��D�^}ʟ\�m@��
1;Luk�
�A�̄�'Z�� K<�1�i��6=�B5AUg���bB�0�"A�02e!X�*ap��4$�\B��������5���t��yIG��D�����.��-;V"<�2Q�l��ϟ��IF���	u��L`V�� 6p���5���I}��'���|ʟ<�����*i�� DP�6������(+�0|�i�\(������F?L>1��O8 ���0��-�P�B<!b�ibVy��C8&@��zE��`�'R剦�MÎ��>��i�8��מ>rx9c�"U7Rrt`�RLa�2�n<*���l�r~ҩW�>l~%�6Rx�	3S��ac-ڛ�|�c�Q:Dؘ�	Wyb�'���'A��'��Z>�Vn��Sj9�!	! ��<�a%�����O �d�O����̦�:`��I���|�6:��D�XV����M���|���
��f���1�4�yR�_}v�5i$H�C��!�F.�y"�صV[���	�y�'_�	ޟ,��>l��e�`��CO�@���b�����џ���Οȕ'�ꓜ?����?�bD�.L��&ϛ�V4X1�S��'I��=/�m�r�&��Q��2.�zm�q�ʲ?�l,��fg����5m� ����m���'��$�R������'�R��fD]�%�н`B/�>�V��2�' ��'���'��>��I<	zNLj�O3�"���#�*����I���d�<�4�i��O�.�:��a�*�*�,d�d�ش��� ����LX�Kٝ9��Ԣ«-	��k<N�0:���e��&�8�'��'���'Vb�'���;�f��~d���'R�)�fX����O��D�O��$7�i�O.��/1,kN"��0V����]}r�'�2�|���LNv�V�P���!�v��ǆ8��5�ul	��D�k&"!K��r�O&˓\bD�zFm^�m`BqA����,����?9���?A��|Z,OҀ�'���2(]��*����+Կ�y¥r�@����O����Oh�D֪鈩2���.�]��$�e� !��l{�z�t�Y�*矒�>��=� ������a��Q�|P0x2D6O���O4���O����O2�?1�.�4q�B�@��|���џ��	���I�O�	�O|qm�_�I�PV�h�Ad�z\4�APME:��$���I۟擫A���m}~B#�#�l�� ��;VE�!��d3}����ݟ�cE�|�Y���Ɵ�����e��2H��p��-�2�t��"�ʟ|�IMy�m�>����?1����_�B��Y�V��P$y c�͓Ms�������O<�:�4������RD��x�
?$yH4! n��Z�f��Dd�Z�"�r��������BI�ɱ��e85)��]��98a�?qRI�	̟���ܟ��)�VyR(mӸ	z��O�0z"|�g�;(� ��C?O���OJ�o�@��c��	�*��t�t�Q`*��q��;4�]��L�	:g�(�o��<Y��M���@���1�'�n�(�(P8*�\�ٲ_�@^�	�'���D�I���I�����P��l�4l¸R�㚘*��#@`�u����?���?yN~�3:��w�6��p�;:���Ɋ�}۞ �u�'g"�|�O�2�'Ed�ˆ�i���ڨJ��U����4JH�\!����'ܪ�UnS۟ zW�|r^���̘�n'~x��d�.
�8�/�˟\�������FyR��>9��?���� M�g�� E�Z�Q�0�+�I6����D�O���;��Z3���3GΜ;P��W�Q&�ɜ9C{���F�b>5s��'L�T�I�|���Q��^�ROH)E$	#u��I֟���ܟP�Ix�O��m] u�v��6D�H9ְC�m��h�>����?���i��O󮉟"�&�8��-�&���h�9��d̦��4��f�"]h�&:Oz�$��
�I�?=a�K1n�=��f9��13S���c��'�������ן����4���W�@1b���$39�|�%&UwV��'�\ꓶ?md��d3�)�O�%X�`C#��d�QՇE �z�By��'��|�'����R��Ag)<�^X8�F���`���"
tB)�+OX�;�c��?Y�,/�ĸ<yj�����7Yz$,[֮�&�?a���?���?�'��$�L}��'�J�B�@�%Y-�T"!�	�b�H̘�'g�6�$�I��DPӦ�+��M���·H(PːlE�9�<iJd�E1&�a�t�G�0 ����<P�H~���ʠIAbm_�Y���1�	v:L$ϓ�?���?!���?	����O��!Jwg��te03��Q�X��'q��'�h��|���1���|rѹ+��V��?�]A*P�U�O���O�FS�Rݛ��T@�- p�T��F낵e�T;%iA��"=��'�.|'�(�'�"�'���'���p�����IE.�*z�xq�'�bP�`��OT˓�?�(�,��#��X�м�5�#8�ڑ��(p�O���n��%��'>A�<�R+H�i���.X�rK(��͓4��ԁ��*��4��P���k�6�O�H�h�~���:��۠! }�ת�O����O����O1��˓Z�&A	YhLujZ8[�
�S�FZ�y��'�2�p���D+�O�!m�R�T�%E�e�4�����(G�h���M��L:�M�O������3���l�<	� ݱ	�@�僟	��]��m��<�(O$���O�$�O����O��'��5(�DW�Vzqz�[�HS&]�\���	�h�IL��̓����1�);��X)�d�	�3ae_:.�fa�O�O1����Ѫa��IQ;��;��Û��v�ۥ`�@%�'�Ι� �D��t
V�|RV�P�Iџ,��ޢ�lZEk�4:T�v��ʟ��	���	}yn�>���?	�C�P��;|=��y�+{R���I�>��i�x��7��[�UE��Z��U-4�-�&���^H���ZR,�� �W�LX'?���'�L|��/by�taf�9c� ���ʘ"��	ڟ��Iϟ���b�O��@�%��Q�qOY�'X!� *��j}B�'��fcӼ��]6$��$B��)j5���&�I⟜�Iџ��tK���'D2T��&�?mB���1ň�g�6C>|����&k�'A�i>Q��ԟ@�	���	</�z�Ye@�=����ƣ'���'0d��?!���?�K~��Da#��F�~(I� ��7
���Z�<��ݟ�%�b>i��c�Ƚз��.`N\�/��q����O1?�Y E��$�"����Z�Jv�`�qF/z:��n�"yڈ��O
���Ol�4���'������X�a��;L�7���=��Y�d�͟б�4��'�ꓡ?A���?1Fh�SE�Z��Y=�8�!`�5���Bܴ�y��'j�9����?I�O������&B˨J�1�D� K�ʥ+G;O����O���Ot�$�O��?]p �E�fI@��
$l#|�e�Dy��'� �S�'uӤ�OH��4cT�0h�]��]>(EԈ�e�$���O��4���x �z�`����X��G��v�Y�+�vl`�2yt��`��y2�'�2�'��	C�E>:-xX+1xY� ��\�B�'��,��$�O����O�˧d	*�kH�3Cޝ�O��+4A�'�꓋?i����S�T�Q%�P��uN
��P1�M�GtU#�@�[֛V�<ͧ�8�Ij��=6b�9(A�(dɒ�ᇀ��PF���͟���ş8�)�KyR�d�8���L$K#*}��A�;3p^`4O����O�oZJ�7��	���z`k�~Y|�p�M�	��@��-E�����*�TlA~"�__&�`�f�� X�"v��J��%�"�	f���!2Oʓ�?��?Y���?����)�֘h�\���+�e��ifq�'���''����'I�7=���
tA�8�� �)Cwʭ����OP��/�4�~�d�O�P���z��4�Xd��O��A ΍�	�^�	�~�L���'���$�H���4�'��m&	i0�`�  ��-B��'��'�X�0��O"�$�ON���-F>h#�)$.��͑5��#���0r�O��$�O��O�X��#��L���Rdi/u(�H3Ė������$��m� ��'I��Iߟ�O�f�؉��� bs�D��P��͟��	���F�D�'��䋠)�1> >��Cg�^���$�'�2듸?��fI���4�}�R�E1W�,�5�Ձ"e� 0a1O^�D�O��I�*�7me�X����LI ҟ�ؑ��d]��� LX-U��q /�d�<���?Y���?!���?A!(D�P�ɍ�E�1a� ÷���t}��'"�'/�O��+}5�,ڡ%N�R�8ŅM�n8~��?����S�'@��[���5>*NiAp�=a�M�� ū�M�EW�K�l�,��/���<i0¥g3d���.�4���g��$�?���?Y��?�'��$U}��'X^���g�iG,�E+�)��Қ'�6�)�	�����OP��O���CS(D�>t�3A��@�2KM�oZ7m9?Y�"̬=���I0���1�1�J^ct����5���j��h�0����`������@y�����@8��a!ą�^t��ba�A����'NBö>ͧ�?�i6�'����P�B!,�2!"���:�B�{!�|��'+�Ow����i���:2�*ă�"��0����G&�c�ra��e��8("^�y�OS��'��%N�B��=["��u�~��K��&iR�'��I>��$�O���Oz�'4:q�� 
��y�0-P�X	�U�'vF듨?A�'Љ��I�2U�tr�-��J�u����7�2H����"�"
����|��b�O<K>9ЂIh����ìα$�A2���?��?q���?�|�(O��mZi%Ri����4C��T�&�ן�	��M3�b�>��:���nǛy��G�U5S}�q�'��B;k؛���py�M>x��T��ky�|L�e�7g��(+�ʴ5h�����O����O��O����|R�F���X���V�~��Ԫf$tS�Ioy��'��nmz��pO�.L�e���9�JIS����M+ŵi[8O1��$A�loӴ�ɂ_
i[F�R�LqpV��!KT扷e�m9��' ��%�h�'r�'e����ʲ$��D�"&Ԝ�C�'�R�'�BQ���O�d�O��$�g�� �AE�p(�iVB�	|r� ;�O��D�O,�O5�"D��b���F�~H)`�>O.���<h�TB� v��'����[?a���H�DDФ1����	��a��?a��?���h��d̝*ۦI��L��Qe��y%��*Fb����F}��'��n�"��s�h�0B�2���D���oy��	�0�Iٟz��ɦi�'d0����[_Z�IQ:�B���ݏ
�� (A�9����d�O���O��d�O��ă ��h
c�ϰ";�UI��J?���Iҟ,��۟�%?!�I�(r �ҋ�J�l�z�$�<��]r�O�\nڼ�?qI<�|�!��'�Hpz��D���� �/XD�i����d_$P�l��O��C�ĉFjH5T��},p�q1!X��?y���?Q���?�'��z}"�'9
yI5��2 �@��*(�:Z�'��6� �	����˦�����MCq�Z��č�g��n��g�˗	��� ٴ�y��'ӌU�C��?��_�\�S���Sf5aP�j���=t���nn��������	۟��	ڟ��*���c��ͻ���[_Y����?��?�wQ��'�Z6�>�$G�y��("�͊Z��a qD�J�r�$�d��Ο�IL/P�\6M<?ّ"ٮY�Z�@+�3�@|	 �@!����u��OF�xK>�-O����O����O�����3���ु#	_j�����O����<-��Iܟd������OT���N�R���g�+*'*�x�O`D�'G.6����%��'%S<7#Ő)2L(J��B�x�� r2�!H�P� #���4�a:��ГOj�q���{�0�v�O#��R�e�O����O2���O1�Tʓ{<�ΜF�V�ñ
��� IP��yBZ��ڴ��'���P�f��*=U�AW��9���gE�DgL6-��m�O�զ]��?��:f*.��_>��L1<(�gR�,\���Ŏ�+}�<Q���?���?	���?q+�Rp���d=�D��3^?H)b�ge}��'��'*�Oblq��nXDm�9jE*�O.ܡ���cF�D�OV�O���O��T�orj7�a���7�؆I�漊af��"�I�oi�h�m�.b�$/�d�<���?	�� ��� J�2蚬�à�5�?�����ߟ�'X���?1��?����}��c�`�x��� ����'���?a���|�2Ռ�����3a�0ϓ�?��@V����3ܴW/���?�P'�OL�d���*���拏,`jaL[�@�D���O����O��d!�'�?��ӈ��*GS�+"��ځ ��?��]�H�'��7m/�i����S�dt��"IDOŘ�r��e����ޟL�I�Y�mZ|~"�S!f��=�g�? ��م.ݞ:g@����:U�l9�W�;���<���?����?��?Y�ՏI�  ��ƊA��13A���NF}"�'=��'2�O>��ٽF�L8ꠣH�窩U
ȣy���mD�v��O�O1�,�*���$	���fD�e.x)����"N�L�H�<��D:~��DB�����D��|P���U%��
��H�!F|�$�O��d�O��4��ʓ@���˟���*P]}�͚^#0�]*�JV��cw�d�tѭO����O\�ğ���ɸ�+�b,dL��M��P�w��=O�$D�"��M��O!�	�?��]*,��M�Xh5�u�[5�T�#=O��$�O����O$�$�O�?����U*�����Z�g�J��"���<��ٟl8�O^��v�|"���N��i�cåM�:x�$�ӘZ��'�r�'��ؐvs�V?O�dX-��PZ����rBֹ ��Įj��cǊN��~"�|RW����̟��	؟|���)q�6��B� �m�'F�����Qy���>���?a���Ձj�p�!3�z���K��I�����O��D'��?��?3��BV'�R�d4c�.M P��IYG�
��}�+O�:�~җ|�` `��lH�fG7��x���3W��'5�'��TY� Y޴!�Tɋw ύ2��5��F jT,͓�?1��]ɛ&�$ry�i�)��ͭY_z��p
M1AW|�����O�6��t�7�=?q���,#���I�����(z�4|����[�� �!��$�<9��?���?��?y,��)�LG.��XSw*�'�0��oB}��'�B�'���yҡa���Wc��:�H�i��I���[�l�йmZ��?�J<�'�"��y"���4�y2��y0���.:]4ͣ�a�7�y���.y"��	?J�'x�	ğT���s|�qFR�Z��ܡ̈́�>@4A�	֟l�IП|�'��?���?���ʤy�dfcH�/���$NC!��'����?����$�����^.!�(��ԋ���'C`Q9uƆW��(����~��'�(=��:*xF�i�� �*�P�'h��'�"�'��>]�I6:L9��K1tu�߻C� I����$�O��dW˦1�?�;=j^X7�n�Z9�v"��f�Γ�?Q�x&�Viۇ7��?Ox�d��iF�����V)ytI�&�<��C�6N^����@4�D�<��?Y��?9���?ل� w�X`S��)J��q� A���Ip}��'�R�' �O���X�K���)�ĉ�<����ӕt����?��'����O+��ش��0.�RM68P���.�3u:p�Q�Hy�c�8I���E��yy���!�-����A������'���'��O��
����O���c��M�L	��N#����+�Om�k��v@���M�2�'��%W�Eٴ��&�"��x �/�)h00f�i��$�O�16�����M�<A������`^�hMx)�ڏ
8�L�GA�<���?����?����?��T��	Y�P�����j����L��'��>�'�?��i��'c�L�w��?d�MP�02�䡉4&-���%�ߴ��S�#�M#�'�M�|�4����5N������(1ZP8��-C�t�d�|�]���	������pq��D�|x� �\�B�T)q�Gٟ���Ay��>i���?����F$)+`](fB@=�t4B��
+�	���ʦՂ�4Y����D*BJa�C"ޟ �����*��R&B��$Č�Na@�!���<�'=M4�$����I$D�񓪅��1`AE%f���y���?9��?��Ş��ۦq3!�9J�������F;,��`m���',7�%�������O�Qy ��XLx�A�/�&e���HT&�O�D����6�}�t�I-t���(��O��E���pҦP�u�L� 	��z�����O.���O����O �ħ|�o���|����@F����6��	̟��՟%?�	��Mϻ=ǒ�C���jI'HJ��&L���?�N>�|�h��M�'N"�����"~@���$�	Ϣ�8�'���⧤�Ο�`�|�T��՟���E�L�����\_xkei�����I��P��|y�"�>�*O����o��,ѐR�#�9a�J�� >8� �,O���O�O���ת��@(8@��L�b��3O4�D
�������(_Q���J+�OhE���U�� ��y��$3Ѐ�70�X����?q��?����h�R��4'��h �(C��������9:���T}��'B/z�\�� w,��P�\�4�@K�;Y@�I��M+#�'꛶@\�-W�����P�C��[O����rq*t�a�*�"#b�5��5$��'��'�b�'+��'{�X)�@ͦT.��[o��M����V���O����O��$���Ot|�r�4i��c��Y�fc�x���gyR�'8�|J~
u�.`y��s'��s���`\�N	��'�#��d�DLn�j��m�ޓOd˓X��h3Bݾ``��91�m��8��?����?y��|�)Ofl�'������r4o_ vd����e��!H�'j���h��OHo�?)ߴ\�n�1�ʡ���c"%��1v�0PQ��MK�O:��c֠��r�&�����|p�S)wY:�Pƈ�
o�EJ$<O<�$�OV�$�O��D�Ot�?�s�+:Q����+�a| �8����������Y�O�ӧ�MSK>�%�\:������dD��f��-~Q�'Er�2�N�MC�O�A�� ހ��N�Ox�Mc�G�O�T��̸�?���9���<q��?y���?�����rc�԰90ΩC��&�?����D	`}b�'(��'�Ӭ�~qPP�57�|�[E(�s�`�Zo���M���'���IQ	=��0����$�o�&"���w�H>��HJ��<ͧ/l��Ą.�� ������\9g��h��3��O՟8���t���b>��'B�7��8�� ���#�NM3хX����O��ę���?a5]���4�l�9�C}��1���T�͞`�6�'-�6ǈ�B��v���hQ)�8\���*OOy��A�)JQ�f��m���٣IŤ�y�T�H�	����	��	埰�Ow�Q0F�K�"�⠃�#޺A)>�WC�>���?)�����<Y��ywσ�d�D�f�����)&hw>6m�Ȧ�iM<�|���� �M�',B��k�*#��%Q�H���"�)�'���0rk�ӟX`�|2[����ڟ�a�g��F���G�/�Re�o\ӟp�Iğ��IJy⥯>���?	��
���s,��t�\��`��#H�<�"Ͽ<1��M�@�x�R���x�Ff�)@A����L���:�^�s�g8����j�K��:���dz�ӉB�%��P;�%��#a�h@��O��$�O�D�O�}�;XwJi�g�2I�Nt��%ǕJ�~0��]N��vy"�n�`���% �����0H9 �3��������Dn�<�?9���'��#���?�;"hܒ-����g�h�@�sQ�'U��'��	⟰��՟��	͟t�	6#������ɽڠ�3�E?Z�p�'����?����?���df�}���ӢÐ�P=����=4��?�����Ş@�$���S=a��iNK�j�ؠX�O��M�!W�P+���~>�d/��<9���1���aN��k�k��?����?	��?�'��do}"�'�����1"���g@�[��z�'ђ7m$��,����O��4�.U)���u_�m��M �u�t�$�\=�7-&?I�)��ATB�z����7J� ��;怙1K+%��g���ퟘ��Ɵ��	����ʃSI
U #"O)P������?9��?9]�����4��B�Pmz5'���8�Hc/܁���9L>I���?�'[8�)۴���P)t�d��W�(z����{̩e��~B�|bZ��������I���"p�V4{3��-�? ���z�����(��~y��>q���?������X�6�p'��&�=3"I��<�ɦ��D�ঝ�����S�d�͞U�ƀ��`�/Ud4a�� T�YU�ǋp�	��U�擒%�$U�	>��9���-cQ\	CLW�`��=�	ҟ���۟(�)�Uy��fӈt��
20 �"��U"0�(��D�O��$�-�?WY���޴-h����8*oN}*��_ n���ۡ�'���M�bg�������O�6��T/uy�KG�eS�=�HԼ}w0��yrU���I �IП��	؟��O3�yHP���sp���%߫[ �g�>���?�����<٣��y���"�b�ӓ�W�@TP�XUD�$v_�7�̦-�M<�'�*��;�E3�4�y�Y?$޶� =]䠸T䒦�y�mۗk6L�I�KN�'��ӟt�I.4�pehӢ	|�H���b��%�Iߟ��	ğ䔧�\�H�	Ο�I�w�����O�2M���M�)����? U����4*d�Fo0��V�fJ�R���-b�P� ��O���>>�ĨCf�ɺ���&?�[�'������&\d\���B�� ���Z>Wʎ��ߟ��������{�O��é!Ķ�+Ѧ��dk
�9FE�.%h�>I+O�dl�a�Ӽ�s�kj>�`$�M-s�$��+�<���i��7�Cܦ} ��ŦA��@-Y�_��χ8x����G�Tu�䱷�֝a��'���'���'���'_��'��M����R�h�h�C�T}vA:�[���O����ON��7�9O��`���7�x�'�m;�X��'�L6-�ԦQCK<�|���
06?l�[dCיy�~��e
�{{`�S�c���D�)U<���[��O��Z�,u:��M8gtQ��L�6�&����?A��?Q��|�*O�'�R)Q�D+��BC��
\���Ѱx�R�y�⟜x�Ox�$�O&��ڮ��`��\�W�f�FPEUs�m��U���?�'?]�];����VE�(�:����)ft�Iɟ�����x��ş���f�'c��Xa-�=p����M3u��q���?a�>��i>-����M�K>Y��	�� b��?~�FaA�吂���?A��|Z��ހ�M��OT����-8�zD)Cm�dUʝ�a��R��բ�'�'���Ɵ(�����[����G�@��@,x�ݘp�'��X���OP�$�O���|B�ʋ.~��Uj7�Uy�.���W[~�H�<	���M�W�|*�|�rp�W-G��!ʹ;�؁�D�/J���pO��0����|�"�O�8�J>yuB�=��acfY"FW|�q(���?	��?���?�|
-O�=l�s%䐫��O4��MA:cIz�yy�g`���|�Oh�o��	
��cqcK5ռ}��HG�P��ԑشb.�V���I
ET���O�h�e�	�z��<)#����P�86u�d���<�(O��D�O����O`�D�O�˧*��ʖ�޵&�zE%��5S��� ]�<�I� ��U�s������c0i����uFm�Qp�����C���ӀY'�b>E�jX���S�? ���^=�NT ��Z!+$l��6O��#uJ���?�r #�$�<���?�s�ܿb���Cb���K�G�?��?�����Tk}B�'aR�'��Cwf�7q�(�AՌ��z�B	zr�dh}r.fӸX��A≰�:q�[)^�m�$n�\7��P�2<�@�5x�p�PN~��On��+6�Hg�֯o�@,jc�E4
(����?���?����h����(rͤ�˴*��[z���FIdk��Di}��'H�jt� ��Z�(�3�_�D� ��cIu��扚�M��i�7M��_QF6�e�T���k ��H��OP�h��Զ]��`�U K#)���3�+�t�	by"�'���'���'�R�6nt��+<�
<@6e�)�剀���<������?9ӥ�c��u�3�ԛ�LI�Bj��\���|̓���|B���!�F����2E�&J
� !�"��Ux�H"�7��Ę��`X���2�N�OjʓT����#���8Ą(�$��g�h�(��?����?y��|�*O& �'���N#,��x��!ɘ�ޜ2�ɀ��y�Ho�8⟰۫O�mڮ�?��4#����6؇v�\C�@�+�z�8��� �M��O�h:D�I �R��<����d�����#�Za �,�H/zY��8O��D�O*�D�O��d�O"�?Y����K���2ց��"dY�F�ԟ��	韌 �O���O�oI�I�q�>��� �=� M��-D��%�L�����Ӫ��o�~�g��0�K`�%s�H��
A�f<�*�)|?qM>�,O^���O^�$�O0(��� ��}�6��Zj=��"�OZ�D�<�wT���	�$�Il�4���e��&rl0��ŋ����V}­l�Fpm����S�t���}A4x�4S'Q�|�+Ӹ���"�%{0ab�X��SU�҉�a�I �P�Ä�+\.����T�F��	�X�	����)�gy2jӺ�;�$�+kF��&�ǀP��с;O�ʓ(���d�@}�|�j�`R'��J�$-ψ=��%���Ȧ�QݴvP�Z�4��䏪_�v��'?���us����5�*P�rFϯ�N ͓����O<�d�O��D�O����|��DΌq���r�ڱתQ�oO��ԟ��	��%?牿�M�;B�$U�� o<c!gZ$8�Q �i 6��E�i>u���|��d����͓
��B`�1a���&#�&!3v��)���OxiJJ>�.O���O��(a�Ͼ���J1�Ϟ�@@+��Od���Ob��<�3[���Iş��ɈD�\| a�G/���p��8;�F��?	tW�|	ٴ6=x��G�;��	Ic��"Pd���>���T3X����2y(j���I�|(x���?oJp2r�!;�d�i2�N�a	��d�OF���O��$-��3 %ͻ���.%V��Ŵ.��)�I���į<!�iS�O�3��hHC$B�6	G!3�����@n���M�⢛��M+�O�<��cS�����q �$�EKQ�Jݺ �Fa> �j�O���?A��?����?���t���/� NRx��C��`�/O��'2�'.��'^�IZB��2Lmp�� �1�Ȍ�ţ�>i��?�L>ͧ�?��P2�ч�
<wN	�G�@-b����T�\&�M�d^���c�:�������%#�b�@�ϙ�����'�4}����O��O��4���}	����<@tFߏ7]�̡gmP�X��x#��m�Dq۴��'3���?����?�4f�B���P"H�t�r��b�B�f2M��4��D��+]�9�O�O��-�8�H��*�q�P(9�y��'Mr�'���'����^>-��#&I��:��vA�l�����O���Ix}�O��wӚ�O���]8D�BCI�	8u��<wI�Ot�l��?���aK�ho�~~�$�?0gN�h�i�Y.�}�#�26��	��B̟0�u�|�W���	���	ӟ$�1�I�#��BA� ΚP ������I{yb��>Y���?����iW��b���K�EN�x{4d�(��	���dIΦm�����S�ą">9��c7��/f��@bogXX �#c��}z����V��9��Y�I�w��d����H��<��i��z)�	��p�Iן�)�Gy��t�NHj�O2�� l,-���;O��D�O��n�a���ɑ�M�c"U"^rX�m � Ր	R3ݨ'�i�"�ٶ�i����/,e���O���'�� ��qBT��4�Н�ß'�����ퟴ�IٟL�	M���Pk�j�O�W�ΩZ��Sܞ��?����?����s����D:4��F�6�B�@&&I�D�Od�O1��i��#g�N�	_�<E�5I(�<��,AG}��	$a�����OؒO�˓�?���S�l�Y�%;H6<�0M��&�1��?����?�+O�A�'���'��A.GV��vL((f4�r-[/*�Ofa�'�r�'n�'�v@�0� D�:�@$f�����O�̑uF޵A�.��Q�)���?�QC�OVR�L�(h���݀{��РEa�O.���OT��Oܢ}B��7��y�D�ԯ%����lT8h}\A��o���vy�@qӼ��]��e���<��P'^�6Z��I��M��id*6m��a� 6�=?S�]�yn���_��
u����O��$[�/��5<�UH>q-O���O����OX��O*tC#+���A�P�%U��S�-�<ɅU���ԟH���s���7l�E��d�pʔD.�iA�Z3��$�ƦiI����Ş'Vrh� 
�� �h�j�s�#	����n=	^�ʓyPL���O0x�J>1(OP!�$̘#z�0ѧ�S !ҶY���O.���Op�D�O�ɨ<ї\���I%[��,��^81J\��B��|]���M[���>iѿi8X��v�>�դY(0Z�m(�����D�C*� qd7�&?I��
�v�I���'���%��x-J%Æ2q�RK��
�<����?����?1��?����)V�V#�٩&��X���ui�'�r�'�2˨>�O�X7�6��1��ke���rA����I�B�Or���O�#{��6�9?q��QǢ�0`�\���C��O*h��e����$�ܖ'-��'�R�'om"��þb�sd��%'�4��W�'k�]�(��O����O4���|��NBB�ĩh�Ɉ� �}~���>���?�L>�O妵��e�u�|�a�@���FnZ�y���Եi�2��|Z'ȭ�@$�P;�O��"\6T8e�N�o6��� ��L��ӟL����b>͔'��7�?)���p�J5���aUf�H��Ŀ<��iO�O���'� ŋ'D<�� 0G"��RҪT	���'��i$����� @�O��5[޸��oX!Ը���&t:$̓���O��d�O�D�O����|� �W-�l����a��} �
փ,��������`$?牸�MϻdZd�#�I����c�[��xdJ��i$���3��I]>7�~���7@̾@��e�壐�."���'v��4�})���\�O�˓�?��S�(��'dT�5�&��ש
 �-s��?��?�*OD)�'���'�"�Cn�><�!=�6�9�%�(@�Ox@�'U<6-J��d$�h����Q�@��(Z�,��s�>?!���:q���&��'�$�䚦�?�q��2W�V�`@n�2�,�o��?9��?����?���	�O��?"���kM�2%������O4��'o��'H6M2�i�%ҡ)�� ���XE ��5�2l�6�a���41���i3�!�°i����4'2���O��Y(�:�r��	�N�XiB��G�IBy��'!�'.b�'9rBUzA^Q��i�"����c��?q�I���D�O��D�O6���$�x���uC�`��ݸG�'@��4�'z�6Y͟x&�b>U�C"#i���Lƿ_y$�iÌ�^��80b��my§Vra�I��'�I*�)k��
E�z��HK֚���������4�i>)�'����?q��D�t�ʄ���Nڅ�ʂ�<4�i��O�	�']�6��0lZ=�ֽYa��6gԂ�I׬ڡDW�1҅�����'�}��n�?��0��d�w@Y�)X�� ���5tw�3�'��'�b�']�'��֥�T�z���˓I� �Q�O ���O�9�'��7�M�N>a5AШy	VŪ�ԓ>�X�'��"V�'�x6�؟�I�8$�:6-$?A5A�("x��g�T!��H��B.4������O 0	M>�*O@��O����O�Ŭ�[���y�/ً?�̊q�̡�?����d�[}"�'�B�'9��I H N�<)�V��5II� ͪ�HS�I�M#�'B����W&{7�]����6m)��9�ve�sc� �|-�Qg�<�' ���F��;��J��L�;�6yU�7�� ��?	��?��S�'��F�=�S(Uh�n�S'���i���S@�p���'̤7-?�������O���@�G���6��fm�	��O�dҫ>�7m ?I�d�q���8��'�^ЪTr��D6�����k��y"]�������������埘�O�x	�f���uNv� �e
�*��C���>-�M���?�M~��$ޛ�w�l(���Q�q���0���'�Ґ|��$�Y�62��9O ��&���N��%kf�P3C)"�q 4O(�JE�x#�(D��qy�O��Dّ$Ȳ�0F@��}N\1��Q�Q��'��'�	���d�O(���O:U(r�
`���r!�H�&�3��-����O��$7��I�`��b�<CR���\i��>y���F��b>��U�'�d��0j�l!8��H�7J�*�l\VA8��	ʟ��I���x�O�R�	�+f�&$.}!D`��,�4f�>��?��ii�O�"Q��u���;$간���Ǎd�D�O���Oy`&fӀ�(!��a���P�RU�?�$�����\�RMB�����4��$�O�D�O&�
8s�UQe�0G� �v��/f��ʓ���ߟ�������J�(Z�9�����D�X�K�=A��B�O��$�O��O1�v�ఁȪ�fm��^3/%�����B�g����@��0	Âh�r��l�F~¦ù�T$��G�>'������?����?����?ͧ��$w}�'D6���+�%���)��ee�CT�'�P7 �	���d�O����O�i���
�����`���U�H�.D�7M:?YW��#`p�I �S��)+WaJ.�ZM�s�?J��3t�p���Iٟt����������r��T&�L�b O��:��RH��?Q��?\�8�'26�,����:\RS��С~�AVJ�
e]�O�D�O��ɡX*6M9?10.�]PJ��#��1t�x���Q��5�%�O�#H>�-O�	�O �d�O�B��I0RJ�� Ʌ�'�� �u�O����<Y�X���������[�T��fB���,n a���ދ��$�m}��'��|ʟ� LY��e�T���Ĝ	�B-CR�Y�Y��DR�~O�i>���'���$�4ɠ&S�*i!�Ȁ�����dݟ���؟|�I�b>�'�6���z\���Z�rU��8ʰ2��<�iQ�O���'��ȗ��x�!r&d�fᐪj��'�ܐ�G�i��I�D�9� �O0�'h���gE ���Y�i��	  ϓ��D�O����Ob�d�OL�Ħ|R`bH�Y�F� 0&Z�A�Nu@!�,$n�	����ȟ8$?牒�M�;o]�h[p�V�Z�1A�,ߍ f�l���i��+��)ր(-�7�~���ß!e��[�.�Q�̪f
s�b�n_:�⥉n�zy��'
�����Q��C�;]�}�ƃ�;F�2�'��'�I0����O4���O�3���0�f��GԠ<,{��,�	���ŦM�����oV����(3�VɹB���u�'bP���kʳ�\��e���
🬛��'JZ�F���Uv��H�9����a�'���'���'m�>=�ɅIN b� �$)�~��%���[rp�I3����O�����)�?�;�����$��'D�x1�cϐx������?9��M�����M��O��7�)��h t��(
#��3gB#tܒO�ʓ�?a��?����?�7��  �r&H=Z��G�y��h*OL��'���'R����'�6�H�,>̒��`Z��D�vN�>a��iz�*��)B<p�j��]�i�^-��@A�� R��U+1���h�ZҨ�O��zO>A*O��#���Al�yi�aJ6���K��O���O>���O��<�Y���I�a����b.	&j���P7۶�	7�M#��+�<���?	޴����c�^X`B�2@��`s�!U��M��O�"��A�"�G"���H�%HxH#��>pNp��2<O����O����O��D�O@�?�4��̚�����d��d�ϟ��	̟���Opʓ,1���|��5 ��ٳh��g�f<jQbڻQ��O��lZ1�?�a�LlZh~R�� ��S#�[�l@=�e�[!l�X�4���8�Q�|rY���	����I����#%0�{�!ؔUX��J����	ayR/�>q-O����|��$G� �\���
	.ڌụ+�<Q��d����4m��S�D-�8(JG䙲?�ԕ�v�Б0�P�ӒkȠLݞ=�@Y���( ��,�g�I�3����,�A��P��lX�'qJX��ȟ$����D�)�myr�eӴ��#�Ҙ[�*y��\�"_Px�R8O(���Op!l�J�	埬K�O��l�8 t�̻�DY�:zDk��G?�	شx՛�`��/K���ԫFM�(;����}yR�̏ƈ�*��I�������yr\���ϟ��������ɟx�OĬ�zr�� ~i��9P�cz��K`ȳ>a��?���䧧?IQ��yǏ�;���{ Nz"�mX2FK�"�'�ɧ�O�����i��N|��@efC������<m��Dtf��'�'�IǟH�I�5C�UZ����\�\����I.Ij����|��П��'������O0���'ԯ�Еb7J�".@,���G3�$�O���'�|7�-CL<��C�MY𤒦��)LTQ���A~bMկSQ*e�1��
5��ON,y��5�2��^L8I�	 �J����IN�[G��'��'�b�؟�$�X*(�2�A�C�&w�M�sfJ�èO ���O$en�z��՟�_Rf���j@��3��2�z���������0Ae'�;?q�g��o��S�#~�@s G;@�r����6�Q'���'�2�'��'�b�'8P��e �
$� ��įOb3�!�W��C�Ol�D�O��7���O�xB�� �l��U�fL-�F��R��g}�'�|��d�Y�{�0����"Th��I7O4:�@Q�i9�˓=O:y"�!���'���'��R�
�5��rYC�6i��OBɟ ������	���Cy���>�i�
����G�~ ։ t���g2Έ��@+���|2�'�T�p6��jfӢ�o*��34�L������st�D"�ܦ%�'{�}�akG�?�:�����w��QrH�@��!��L�8�˙'�R�'[�'���'M���4DW�!Ж�j ԱI��<�L�Ox��O�=֧���'�h7M<�D�O���]�&�J���iUB�e≝�M;���p!�6�M��O�Qj�nR*X���ШG+��3�m"F�����h�O˓�?���?���Q��蓭ѭu~���l
��OB�ĵ<�$T�����(��w����p�>�;D�ːq֜�h� ���W}*p�@=�IG�)
q��8�p�i�Ȗ#J�xU��AJ���@�D�V�r��,O�iQ��?��2��	�F�TZToͥ8�p�i���{.�d�Of���OF��<i �ivN�iQ���x�\X�CV�h4���'��'Yf7�&�����F�3��j[:l�nؓ��)Ŧ� �?�޴.�@<k�4��ݵi�1��w��T� |"��>�ʬ�BE��ϓ��$�O����O0��O��$�|��A3q��h���Ш	���  ǵ���ݟ@�	Ɵ�%?�I��Mϻc.��G�yj�	Bč�y�`;��iX��-����3Uz7�v��G	�~�'hR5R~vx�y��@���x�g�E��Gyb�'�2�ܩGLZ�[��p� ``Q��%���'�'��I�����O���O\�����	 hJ�B
C%�����%�����ɦ�����S�? L�C�&�@��Q �P�yy��:�����T(��;���k�Ӆ'r��� �5� n��5p1�U�)J�0��C��	՟���؟F�4�'q��S-�V.�uڇ ]&>,����'����?q��	֛6�4��d��ߩU��������FL�������ߟ�oZ ^�o�Q~�%\�A
H��ӌ��
�$M\k�x¦R3�UAP�|�V���Iğ���̟h�	�� sH��2�$hH�����&�cyr*�>���?!����OA@R��8�f�cr�&�aC4��>��i���1��	� Dΰ��v�4=0-W$�?&��@!���hi�˓&��!�Se�O��yO>�+O�	z�Aڙ����C\0pVT;v��O��$�Ot��O�<��X���	�ez`K�D��E��<R3�Ӻ/��I,�Ms�2-�>y��i�h�Dy��iB�&A	;��Q@�F67�t�D�21\7m4?Y�m�}���O3��x��YX�' �H��3$}�D�� ��kf�����+ozPpfȒo1��'%�8	�' i�iQV"��G>Ja�ħ�$R�ܨ  �/Q�$�p!!уE`�=��O�-�H�t� 	.j�`e�٪Iݶx�0��F�~a(�Ԍօͫ{�^���#Լzzd�b�(FqZh�v*j}�fŃ:"�x2���o�f ӲfBA��"nV��m� ���k���:�|��"o�W��$�I�l�Ԝ��J�5�.��J���1�W��&�9��m�C�D"2��B>����AI�vDt���eb���㦍��ӟ���䟐y�O���?9�'�Ҥ��Չ�C;&\�i�}��Q�wi�L�yR�'���'�4]��CA����cI</�<0�7-|�t���O�!�'��	şP'���t�P��%��J1���[|��T��=���!��?���?AO?�&d�)C�Z�)���\ӈ���x�A�'��	���&�H�I���{�ٌ	����`@CLX��!F
�Aw��	E���	�P��ş�'?a �Of����L"c\�d���P�J�a�۴���O,�O�$�O�ɀ�]�9 ޅb��+�5�0�@�.�yr�'��'���p-�O� �KGh@p������D�6I�6��O��O����OV��2`:�I=p��xe�0D���k!$�.s�6��O������d�O0}�O2�'���C�ΰ���+i��$X1o�m�jO�D�O&����6��r�Ġ�&V�Q
a"�j+���T'�ʦ��'+u��	��M����?9���?��_�����V�*��-KЀ]0I�ph'm�2�MC��?�'�S�?QN>.�jL���i��5�'�@�b>�4OO�x64�1ڴ�?�c�i��'m��'������<��U����
����5aF��8�l�le�?1.�]b�>OX��^I�^	rd�Y�T���i���B�Z�n���,��ӟp�I���Ĺ<���~�G��@��T5Ė�(X�=aTM�&��'�� S��'��`�'���'�2/��q��p��,�6��0�9j�F7�O��F}^����J�i��iV�I<t,�� '��\��!ZrI�>A���<	���<���?������8-'n,��G �2�~��g����6�M}�]�D�	s��ş@��?Tr��򒊃�g��C
�~�ȩ�b��T���w�P����T��J����:mB�SƏ)�B�AV�X��M{(ON�(���OL��7X� ���-�$ �6o׬	5P�@��א_��#�'�2�'M�.��j���'�$�C��B�Mµ�M���UwӪ�$,���O��D�Qؐ����I����\����6V���3&�t����OLM)15O��Nz�$�'�"�'���fBY̺)@���:?�d@��g7��O���ܑ\�F����n�qC�$ϲe��1D%ߑN�j�nZ�Wl���� ڴ�?���?��`G��qw�$0f��_�4�"⋣SY�7ͮ<���?�ß��Q>� �c�N�;E��ՈLk���5�$I��i�B�zӮ���OV���O�T'��'R�5)��O)H�:i���v��o��D�	�x%�擘r������j��F6�A;�Eр}F$`�����M����?��?��xʟ���<B2����%*��!�Bg�5��7-�O��O:����!��$�O|���O�dJ�lU�,�0䂀t`��2o��������H<�O�ɧu7��|f�{"��mt`Xc$�ܒ�ē�?0�AF~r�'I��OJ�-� �Яږ*��`(w&]�S|��U�<������?y���~R���+4B�ʐ	�b�j��ߖ�Mˀj��*�̜�'m���dS�h�'7o0�K��+;�E�Ao�s �Ao�����b��?Y,O$���im0\���t�|öO+�8Ł!�<?	��?q�������O�U{��S�J�U���3�1p��y�?�����ϥLv�'�R�0��v!��9[-��	�F��M���?��D���|��?����df�H�.�X��'L�r	;v�Nt����'tV�����!��\|��"QO�����i"]+�[���I���	�|��kyZw�f��g�_�P����"D/���4�?�)O��2��i>]�Äi�rd�Ee��Tj�:F��lS�i�ǰi�rAc���O����O�e$��'!��Ч��{��ٱ6�ngL�n����I��X%��S�D)8�5����K��2�`��F�؃!=���i���'�2�'��)J���C%Y3-�dYB )ՕUp"c�j��O��i���$�O���O�$6k 6	.t�)�ɪ~�:��.¦	�����BM<�O�ɧu��^/d�HM�����H��|IMX2���?Yd�E�<���?�����3� �|JW�U(!ja+���|�@MQ&�i,O��D�O�O��Ӻ�@8Y����U��'у�̦���"	KT��?���*,O"��<}!��³��.+�}X1�ɵ1�V6m�O��3���t�'�1(شdA�D��n��Rx�	�� p���;O���O����Q�5����O�Dc�E��UG��g���a O֦	�	u�	^y�O,r�~J�� p���@��E*3�Q�w'�Φ=�	�L��	�@�ɻ��I�O���Ok,J�?d�t šK�2/��P�Y�`.�'d��L��b�s�֝�{6$�ӂԋbp�h�c��
H�69{��$�Or�oҟ��	˟��I�����fTKTfJ� ��w"0$֔�ɓ�i��'�pу�O���ɐ%f*�nؐ8�>I)˂H#DQc�j�t뛆�'�f7��O���OP��l}�T�$	-YP��A�s���Ua)e���M��T�<����Ĭ|j@œ�|*��'�*�b��X%O:�"��t6e1ӵi "�'�b�'�������O�Ɏo�)�b��-�����ի}B7�<���]��Γr|i͓�?i���?�֨�#M�h�Ӎ(�tZDW�/����'�J�>�*O��d�<������0�J@5B8bg�9���GĦ���K��	�X&��Iş����h�s��X���C�*[В��1�F(�
6-MY}�]�T��^y��'rB�'HZ�3��]e%��hIC���yB� 
.T2�'z�'��DU>��Om:��3F�bT,�1��vE�yܴ��d�O��?A��?�� �a}2��8Z����(�.�T�4��	��d�	����N|��Q?���8Z�V���p>Y� /!.�T��z����<���?�f3��̓�?���B��)�3� :A��XQf�L4�Z�PT�iYR�'4Rhҟ'�R	�~����?���6�Y��A��4e���G��q�@\B[��������I�����d�?W�;Z��� D�4��y�6J�M"���<a��Iޛ6�'J��'����>��sy�\�3o�5պ��AI�M�`�n�ޟ����wJ牍��9O�˧gB0��Lq�\�D��	F�|}�e`�3c2��lП�*ٴ�?Y���?��-&��@y�Z��\�r�ٟ&�<p�!S�,�b6���[��O�����H�����O.�Rl��c�Y;D�z�+��PtH6��O|���O��d�I}b[�d�	~?Q�ӅU���
�KW&l<�b/��m�I[yB�� �y"��4�'�r�'�.��sM�,D8�mQ��j�4�H�jsӬ��O���'��IΟ8�'�Zc!�Rc��0S*\��ƭW�� �O|�2O�@��)�O
���O��d����U��Ǔ�W�$�s׭@Q ��#1�i������O6��?��?Q�OS���S�+dB���U�W���̓v�������?����?��'����|z����fF
���(���ѦY�'32V�\�Iӟ�������a�����"κ|��v��3���`�O��d�O�� κ[.� �OZc�@0X`�<HpP�@�@<����ٴ�?�)O����O��ā	�i>7�S�`�
�r�'��8����~��V�'c�����yB�'),�'�?���?�V��[�ȡNS�3� d��
Z�_��	Ο�����,��b����y�۟\yP!�P�h�=;�,�~+�ك �i��䑜'}re�|���O����O~�ԧu������dD0.�����N��M���?���@�'��S�4P�7mŭ	\x�H� w�΀0f�N"���';7M�O����O��d`}b\���`�^ˬl��.ެO{��pg㎫�M�N�I~�R�0�OL���O��N�� ��G bM�h"['�87��O����O����g}�U�L��K?1�� G����锓E�q��_�a�V��i��Γ�?����?a��"a��	��0�eR�J��!؛6�'�rl�>A*O����<I���5��y#�ɡgW=~�*�F[V}���y��@�%���'^��'����uw�!Y��!��1y�`�h�,�M�T�8�'�X�<��͟@�	�w桫T���wb�,#PG	��Mc��y�l��i���	����I�?)�O;�擛����M\�*���&�d6��<I����O���OI�bT��(ѦʏV�,�!�X�eNeiE�4mlb�'�r�'���[����~
���2��!tp�QU�[�,ٴ��1j�Φ���jy��'�R�':t��O��Ic�(���	O( �dx�Ɔ��6m�O��M�P-��O.\�Of��'��B>GPl!r�+�$,1F�s�Cܷ=����?����?�Zc��7���?p6D�e��ɫ�m\�P´�"'�{Ӛ|3@3O���O��)�Iџ ���ҮO�ь�أ"EԖ9�R�׆��
����'U���yr�|W>�Cp�y��P�c�ĥD_���`χ]�}q��iIZ�6�'=��')2�>�)O�؁�"��@;!�X5O�DPy��Z�y��|���Hy�W>�Pfh>��	`��J�N�
R�e�G���^��۴�?��?1�J{��Jyr�'���$���$�\�d�`⭘�7���'��I�`��牭	��ȟ���П q�%;`�I��%��v��U�� ܛ�Mk��?1�^���'�RY���i�]��B�:МuZ�j�: ���Ƽ>��A�<���?����?	����Ӻ�A�[9 ���pO5M�����L���0�O�˓�?�)O��$�O�DJ>>�4�X�IυOhD�Z N�q0$��=O�si�OV��Ob˧��I�|J���b�F�R#��'3e�䛐�����'�bW���蟴�	����	#;�|@o�*��|�D�-vV��`'^ǟt�I�p�	4�u�'�rC�~���� >i���!��-Cg=9{ft���i��Q���I͟��I��	ݟ��ӺFľodB�Iv+�.gg$M�c�i�R�'7�� �'w��~����?���iTJ�y�$�I�8ђ#҈W3���x��'�RlH��y��|�ӟ���%�Ż^�ܤ�6C޼4�85�a�iA�I��'�R�y����Or�$�O�<�'@����;�p�h�XX.P��4�?���c]h@�������i!}_��D�*_��0�W�2N��y �,�Ms��j��f�'bb�'��b?�d�O^��7��07¼-ȱ$�	ݦaz�H�)J0�x��$�\�O����'��L�$�݁�H��t=�<"�N%/�6��O���OD���]��?1�'��T)bo�z�@�Q��z�4��=NN��U�Γ�?1���?�R䉷,�(1�U=~�6Q@S1K����'FB 9��ON��"��Ƅ����T�D�;!L
�Sbm�f[�0����ɟPc�d���Iן���J�I�q���Dތ+'ņ�#����!��ɟ($����ɟ�B+�-8����Wd��K��Ta���C�\��	��	ԟ������&?*�O���0c�k�4AD*��n�Zt)�O$���OޒO&���O
���T�$[D�I�8����\wɞ騂 ��y��'!��'�� ��O��	�2iЙ	H�.s��IEn�9s�6�O �O��$�O��n�O��'��5sD���F�DT)�dR�a$�H"ߴ�?a��U�d���?)�X?��	˟��I7G��q�U�ݱPV���@\2��N<Q��?I�-�?N>)�O�Z�3DJޔIhx��ME�!���4y�4��?��i�r�'W��'z�E���KaU�L����W�ˋ9�:�n����	4'�x��f�	^�$f��M�@�8�]�F�ؘ��,��]���M���?����?�t��b��� �E�)������ZLh��ܴ��������)�_���O� XTOC�t,�Y�	�J��XA䦕��şD�Iڟ ��}��'���]�H>�3�%G�]��D	��GZ���|�Ý;��F�y��'���5֩�C)��c���R�������MS���?Yu�D�Ot�Ok�A7W���;��͝�D�����	�;h��>w(���p�	˟���Ÿ�%8��[୅�Y�t�H�i��Od�-ړ�~ro���b����j1P�Q��M��6s�MΓ�?����?�L~ʁ=�b�hDoP-{.|Q�I�$ �,�@W�$��B�'
�I֟ȢGM'AP$�	���C1j,�Rd�1H+���ɟ<����x[w����(�Iϟx�d�%f�@�+�d�,]ʼ�E�ϱ�M�����?�/O~���x�-��sO���v�J/C��%rE�Q��M���?� �<�C���П(��ȟ�9��҇g8����%/�<�U�ݤ�M�(O*˓8��(������Y��UX��Q5���:���6�M�ÄG�?����?!���?���?����?��$�W�zZ6ǖ�z
)�c懽@\���'��	�L�"<�'?�dn54F 9eP� �<���?v�6��Onǟ��IݟP�ɝ�ē�?�3B�'nt�yt"[�(y��`$��p��6�C�O��+C���I��q�_�S������>������M����?q��?q��$�Oz�	�#�n� O�	�Ҹ����(ʒc���P�n�x@2}�p��՟��	�[�@$p�i�89F��k�(��	�D��4�?�N�'"�' ɧ5��M�!>�iI����5�H3`�'=&t��'r
�
�'MR�'g~�����<w���I�65��4h�L��UɊ}B�'F�'eR�'�b�`��4OfU"Y8P`����bY��y����y�'��'N�O��蠑{�d4�����$�<)ѶO���+�D�O���I#=L�I�
��2�U�]�fIc ��0�|�P�'Cr�'$�!8��l���'����DX���Ĥ�4� �BT�h�@�d)���OB��X���'���Х�U]w$Y"#�Ż5�X��4�?	�4��H��?�[?��������	]%jxYb�'>�� 4��#Z�E�N<����?�gLL�'��)݇}"	o�+%h>
d��"!�N���y��'��6-�O��D�O��$IP~2�ٽGn��G*	V\+�m��M����?���@���i�?&1�V�!w`9��"D�u�<
�+�M;���?���?a���?�.O�'c,ꕊ���Lp�m���W�B�:V^��yd�<��|zE ��<��-��D�ᧇ�0�$��hZ��|���i�'B�'�O6�'�?���>[4x �(,�x�ґ�ɇXg�OJ���6O��+>O����O2��q����!����\�sea%Mmߟ0��Uy�h�~j����?��� qh�{P5c����1�x2��iǤ��'#R�'��O#��%�֨�d�F�I�
!����>H���'���'���'H�'���OnxKu.#�x�:�X,]8��*�iVP8�kȰ�yr�'��'G�O-���]GLܚ��eM�`�S8f�ꓡ?a�����?i�{B�׬����M���T��0bՒ\;��	��I��2J|RbS?��ɭ޶HC����C�^�r͂X=�޴�?�M>1��?����|�OH����j/YVYHÁ��:Mo�������t���	蟀p�����O��[�Yd@)#F(6�pƈ�".�4'�h�I���,u/�<��4?��R�N��j̘��E�tmBo�//5*��	ݟ���؟����P��Yy��+� �|���+H�<��0C\�k��qQ�i�Y����c3��|����}6�,Q|`%p&�$3*�[ABv�����E��̟��	��ԀM<)�Oo��cfMA�>�L��sH�?^��4O=�������yl��yr�'��
a�Bs��)�oK&<z�\��,v�
�$�O��D�O�˓��i�O��I,\V�!������\j���S��89��d��K��F�<����?9��+�|�@���sfnX���ҕn�B�
�i�r�'��b���In�i�E:)ˆ1�&�sg�9n`�ã��>����<)����<����?������n}��Sp���{�DYqs@צL�7�s쓹?�L>1��?Q�k��-��%�e�/�|�;F� B햀�%	&�Γ�?���?�M~b�>���r�5/|�����$�rt��\�p��ϟd%�t��ϟl�M�>y�>Q�)Ї����,�f�Ixs�$�O ��O`�&>�訟b�$�wאe����\׾A���8!^xinZ��&���	��!��1��
O/����Ȏ��uC��8w�7�O��� ���O�)�O��'��#�79!6�Β�� �aX�����?����?9#��<1O>��O��|���^�W� ���*s4]:ܴp��,��?)u�i���'0�']��Ӻ�(����7(�&���h�DKߦ���ן02u�t%��O�y�۴}�°���vj���C�`ꪴm�֟x��4�?���?����	\y���T雔��K5�u)�_<1�h6MS�!��IPyrU>)� J{>U��D'Z�am��+�BÆ�[@��-�ش�?i���?)��y��iyB�'����96�~)��I�h�H��GӘv��ny�	�y2������'Tr�'m�ї��y{n�I�<:,����Ӱ�d�O���'��ޟ�'�Zc����t�,Yڤ��n!4u>9�O2��7O�\R6O���O��d0��+�7�l�#��ӧW&Dx(4�
9�M��V�\�'�RZ�X��ǟ�	�B�b���ʇ�6(H�%E�" 6���aq��p�l�������E U���18 �^�
�qJ��G�I0���I@6.���b��DTy�b��k���A�e�&[n�R�J�}XnH�NO.N�a�rd�_�@��W�&=���G�8�)�䉖�t�2Î����H���V<u�E�dFD��j�Q���nB���,\?\�Dmࠊ:��`Z��Mtc�����#(�3+4�p��N(h���Pc���
��s�
yx��"&�܇]\�"�,ȪU�"%;QO.��z�@�),ڪ����}�N=Y��P3lv�p3c
E�{���BRh��$Z���'?4a��&�$)
�(��~"� ��'�"OX�:�,���d׉DN�ԧ�i�|"A�!P ���ę8��A�N�V�DC(KW�͂Ǩ�Et�E�䇜�QI�-��)�}�8 36媞����/�O���)�'�?1u坢T{Jx+���<�a�e#Tf�<�#��@��T�T�L4-{����a����D�#1 �CG 8�̓u�H���'a"�'� ��O�'�P����,���
�,Ԣ�B&֦(�ӎ�+��	"����5�$�3���k����I-,��n�"s�ձwG*��dK.M�V����L>�3$�+��4 �C��bev���Շ�?)�O��P����	�x]��ԏ������+ZGnB�I!`�f�E$�?*��DÂBэ!Ed� ����'���+w�X2����
���&�<*Q�}JFËŦQ����L�	|yR�'�23�����Z=l6q[�Ɂ�>NRH2�k;p�vmb1��Q��x� �)<O���򅁃T\���3���N� }�T&�976ƀI4#����G�><OȌI�C��t?�v��vʥa�,�6��'&ў��?���U1j�&X�C���ճ�-�O�<ᇤ4  �Y�ꉬT�j�{%w�+>�	yy��+]T|��?!�Lö~����arT�ӷ拞�?i/O��D�O��:��	pG�E���'X�9[�o�STF����3F��E�Ǔ]9��`�l�8g�Y��O��[����ո#oX86� Ԃ��'uf<[���?)O�,{E��8����0h*<|�P��$|O�ݲ��X+Y�(c�ɇ(r�q�OR m��+�$����:
�,�q�@DH��I[����8��֣
T� 9�v�9���R"OEᄫ0y��i�)4��L�6"O�a˱GQ�t$��cʏGOf8b�"Oj���*MH�u�w'�k�FD�"OԼ9��]� ���y���o�U�4"O���e$=zl��Ú)@��XcP"O<$��A5��yiV#]�}z$(��"O�4*Q Z)efb`��"C:1f~$3�"Op�YeJ��}!Ya��>`O��a"OhpJ6�
a����"�м�U[v"Oܩ���	;�(Q��<
�$�[ "O0]�Q�@�9�R�;� �~覤�A"ORqu�[�>6��k��H�T<I&"O� ����Lڔya�)H��űU����"OHh��D�F*�P�FMc�� w"O� Q��7
Ra�5��{	�ٛ�"O�|PK�'Y]�	0I
�
�L|�"O �UlW9Nz��eh����u"Or���t�N c֤�v�p�"O�`BH�-|�Yʥ.B'����"OH���� t�TpP.	����ڱ"O�哰�pd�(cӌ����A�"O,�PdmN����rb��[��� �"O<qô��)��\[dQ�t�4�)�"O؍@��ʖns�4I1%ø^*�8�"O����Ǚ�k����nìdad��"O��3ԭ� @�X-`ToX�pQb-qG"O 8YR��N9:�@W�`I|-jS"O)R"�x&XPq���L9Ll��"O���b�D6�Ƙ�o�81zlB�"O��Ѵ@ѡu���w$V'Fء�"O`eYPE˽5@r��w_iިbg"O�Mj���#_@��7`)O މY"O���5j���z��Ae���^�bp"O~��c���
�
�QD.U��{�"OLh�E#P�t��CΉC��b�"O��Swn��A��Ls��K�7��@"O��R�AG�["(��E$(-�1p"O��{�m�.z���q5O�KƄ�"O��	�I.�1��@ەm��U�"O"�c���IĂ��pB��]�H�2d"O4MX��B���t�şn}v8hc"Oj�DыS0VHQc��IvB���"O�x(�?FRmw��?uiX��"O��D�H1�<aF@>h`�*b*Onqye��:0oz��$�X�$Sp�j�'�b ��IƱK�vIקO��=b�'}"��8-�AЦ���I,����ē:u(D�d��rr:4�u��11B���@	�yBMϭߪ��t�ÙT��Tö�'}����p�KL�S��?q�-�)y�) ӎץ!yX��	�t�<�&.ͺ1�9	k�\t.��fUv?���H�\��|R"/o6�	�aE�R� �(��٢�p>�D�-c��䙻@0&�K�$�7��ے�ҦN�!���(,���C��[�KMҩh����Q�P�!��*����cC'���9`�կ��"O�p˔EH,�5@d�ǫK����H�@���}���'����	��5]��*�M��QC�̲�'���c -7X�0%��NrJ:�'x��b�!�O�ak��#�$���������'cDhB�����"p�ҼQ�>qk���04�N�T,!D��w��(q)@M�"�_�'?h1kU(5ʓR�B�P���5	'��KU���G9o�zB�I�P�B��5���#�\eP����*�O?�DE3uzfL�w�@�d�l�#�'5z:!�$�����#L0M|�s��чh��d_l�'6�$��{��V9`Y��/<	:�#@��p>��38���Ie�X*3[
�� %`X�8Ҝ�O��@�`9LOĈ+�G@�|(�e�e�2C�8����	Zj�5����'0�]�r�F�V&|Xc��^�`@b
�'���#V/H�I��
j�Qƴ�ۉ��Y�$�6#|Z5�
0M������x����I�<qc�Wʾx��Lǜf�H�#�SOyb�
1{�OQ>ɪ���V#<Xj���C?x��B0D�d`� T�.Ð��HQ���7K-���LY����p�SI��A�\���H�*L@O�Y��i�6De��(��73]8��%��$/�!�� ���T(r�(�� ˝H����S"O�M�'��{����1���8f"O`���恋|���7�ڳ7��;�"O��'ø6B����g�"I
�����'J���t�d]�g.���s��+ھ,@��S9�!�$�8�ò"�	�&m�e�E�1�'�6M�����L�
�j��`�9t�|e#
9NC!�$���SR�V z��h�VM]�,D�O����)OK�BH�ʲ��-(\���K^2��x!A�P�X�ף°DJ�1�E��u�JO�e��Lӄ7�"���b�&���2S�'�2��A���^�X�BA��=��Q	��I�w�!�¢3!��#A4�����J�n�!�dK/�$�� S��#����5�!�D@�7<�r1+��4Ih3���2�!�dՒT~P�4ϛr��ԏ�=�!�d�����kPڌxf���D�G�!�dK=R9��x� �=@GJM2�^#V�!�J�nZ���CV�#B���&ͿC!�d�C@}@�0y�\�!tN�p�!���*�=�䎓u���#S�!��^4T�Du�V��C֐`"��^�!���'TA��)Wǟ�B^��!کi�!���%L���`S�n�҄����\�!��N�H@�R�����(�Z,m�!��ά!ҡ@U-5��TГNL>'�!�$AH> ��&g�E[�*h
�'$�9`��I��L���_���	
�'��B��sx`gd�9Y�<���'�z3v���B�hb�.E6Pxͪ
�'��+�LU��.�[6l�M�,(�	�'�J��S��C 8�!6��1`��Q�'�XM˅b��!�L�"6��wB6d��';ưAu��cD��!6`ω
��'����a��"��u�� �\a��'����GeNzhRR�X$)�*|�'�m���,Q�y���LBI"�'c���$,�\��@ck�~�f3�'M�M�#OY;QX�R�K�n�zh�'�H);�U�!�@/��d�����'�x�P,�������L�JQ;D��+�B�ˑ������<ai�.N�H�*�5�X�"A	WyR#�,�<�"	�J������ �]���Y���'I���ʭ*���j���O�	���i��������n�HN�X��$3\OnIr�)I�	�$�'�&eCS�_�gp��(�H^�}c����°M�����8§G� �;��� D`��x@�A<&q���=aU �<y�2���K�O!8!�R�5L�I�QKB��	p��¦q
7��;-9�')�#}J�ʎ�m�ɫ7j�|�`ݙew��蚦@��~��Ɇ��Ӫ��,'�t*я�)A@n�񱍟�B��\�����cc=a��]��	�PL��#�S�nw�Bd��t������U8�.���� �|YB�a�K�\��'}ם�"M���S����������U��,�m��	��y*=�MyÉ\2G:�X`#�_�%)�����O��%v��X�*?
�m;ǁ<}2<�l�P2h��F7x`�
f��0R�'L��d���X�\�#H�2=���3�[1H�f�F�7y
xcW��{��%�(�F�WR��O��8�X�j�������R�p$�W�	��@���@ |�ecu��&����ѕU+�r�eE?^��"Cn�ly����h���	_�f���J	 ��]*BfR"F�6�ό1rR(#����MH ʘ2��O��p"���n��z-r���(͐'8)D�P�Q�R�O��h���<v�2!i'��_�.��P霶X���a�$�6�<q���S�KqO�N��z�ʓ�LK��*�!��0?�^��	��lK4 ��:7�݀q��(�cN�QN�Eqˎ3���'"�2�����m��
K�%ҡ:���Ԣ9��r���
5۬��jY��?��8T��	�'�* ���g-I��vB�ɒ,���玞I��J��F"`ϒ��ߌ1n�Xr�lʍd�h% �$ٲl#?�� J@z�M���l�dڨI�za8�"O� �e��&��ʵNA�����
��6M��9�(j�ϲPPZ�g�'�,h�h̚L�� sꐖ`hؙz�6&�����ByYK�N�}(�i����A��(�O��t��Ն�I�`b�87�Q�	��ڇ�ӛ
-�"?�6�'��ep`3#H	�����:��A�ȓz�,�cQͥv
�I���[,K���ȓ��(A �-�* x�G�0xe��ȓC!�}����<X�y!ܩ��1�ȓ/�~���A6_p��d��K|��
d88ӦA�p�'hތUu�`��B����6*=�`�Pd�]�fx��'��E��iV������<ꀆ�i��йfD�-8�p,zWJ� �L��( ���UIɏVd*bR��AJN̆�@M�� �XB��T�J�e]4��ȓS-���PN�0��IЃ�
\D�X�ȓ;7�EGÑ�M��`��ǽzx���&�t�h���1�P8 / "z��=Up��/�r�Vb@�b~,��0~�f�J7V�����$r�Єȓ���q��7`�H�{��(�����I����r����sm��ȓ7n�`Xa�֟G�.��R�"�>	�ȓ<�V�P��&��8r����h��ՅȓY^$����в��b�Bжw\���ݺx��D
tIr��@X}�q��|
l3!�J✄��BG�)�ȓKk�D	ɑ	n�R�rE�9fb�ȓS�}A�l@4t�V�4�YR�����F&a!�B����Ҽ6o��� ɠ��&�Կ}�t�q�=d.��ȓ1�1��H��P ǃ��(��l��%d)�Ct>!a�B�qJ~C��1(��79!�P,8ЬC�r��ȓLX��9`*��>#�|�af��U`X�ȓp�����b�.��h���_�	���ȓGh���U/76rI�2"O;a��T����ק"l�x�'ؼWՒ��ȓ^T�(�#�`����wH
��ȓb�(C�ȁ#HCt�ӥ�-�E��E��:��N|���'SǴن��؈��)�0�TK'��2sr�h�ȓ�%17�4�;R�\0ea�|������e�+���2���*'�X�ȓ_n��"ѩm,�B��+u�,ه�='ڡ�u�N3?��y����=b��ȓjj$V-�!K���3$lْ'�-�ȓY<�I��A�9=���a�E��ȓ����u��21gF�0�S ;�L��F��DH�B��k����E�����ȓX#Z�1�K 0�� (.D��ȓn�h�l��!O�9��!�,:��	��/Ɛ�ע4\�"�� �Cgڤ���6����"J ��fΘA!���]�@���iD6�l��2�ռ^��y��f�CV䁣]2܊�+K<��P�ȓ~��GI��?|�T��r��i�ȓ9��L�$��	4�9F��	"�Q��Y��rT�S�
� �񤈜0[�\l��� �¤�2�U��a\"�ȓf���I���]���0���y���<@8X`R�J���Cߴ�y���'g�܅���0=�~	kc#�y
� Ȅ�ܸz�d���� &�$��"OP	�%�#!�&)x���	Q}� "�"Oԥ�a@^U$x3��_a�L	�"O�T�ը�^�]K��D�=}@��"O(�� i�+ �*��T�`4��"OrE��R//4�y2ũ�=��@p�"Oި0 �&[p�7)	4Z��B"O\	+��FZ�(!K���+X�Y˲"OD<s��L�\>L����>��5"Om	Ҩ�#i-Ԕ���(W��R"O�)����?xz�ܡ%@�8�b�[�"O��{QmL1t���8��K�kİ$"OFe	��
z:Y�����Ve� "ONk�H�..��&.��
��T��"O�![�鐧,	T�M�8#DA��"O�Y��=L 
�*7��0
��a�"O��1&M�7&լ�9aD
�X3"O>8�兇��9���Ն'd�q�"O��)��� P8i)C�%!�Dh��"O��'*{nhVi߫r����""O PaACX�eޢQ��O��{�"O.0H���G(<x�5��&I^�Y�"O\MX�\>@"�i)g/Qx�c2"Oh ڂ,C!s��y���]�v\y�"O��! ��Y��X���5]��ab"OL*��2u��E �M=,Vc"O�q�G��q�S�懛XĤ�:"OvQjbM�r�\ �Y=��M�"O=�I�&'����sh���TAse"O��`�YW�� �ƈ"m��{q"O�X�7]\ڴ�h���<b��q"O
`9P�ΜLv����Q3p�`�"OJ�*���'{v䀘1�L?|D@XB"Op��BhJ�gSD�-�4&>�9pF"O�|X� չ H�]����1%FУ�"O�K����i"J�r��\�l�"Ov4�p9E��A©��uV4��"O,�g<!�ݛ֎Y:f��"O&�P�(�mA`鹆L��(����"O��з���*�
����#V4��0F"O\m��G�?3���J!Q���'�y�Z6�x�"$�X2 � ���K/�y� G�`���� ��v�iC#�"�y�� L��U/�=y���9T_��yr*JTLZ �ѦK�vMx�!E���y�A#bCҡq6��]�0�j����0=��«��#�u��N�!W$*����)�y�N�l5r�KՖ/v��A�yr/��Z��K1n�7��u��$݆�yB�2`�傡�.
6ػ6��y�f11݄]�uB�mVʠ��` ��y�������7-��l�&@&I��yr�A�y��H�P�1)*�
�&���y����u0�yFh�8rV�0A��C�y��
|7B%1��q
u����=�yBdK�N7,�b�ǋ�c憤p��8�y$Y ����!b{�8�X��y��L��@���_�Rc.T�v%/D�<ADG�eg��+�璁6� {@�'D�䀦@dy(�S�*�>�0!W�$D�j��@�42d� C]����<D� +�á��|���ȧ!���"�g<D��H�%��u�rԂ<���0D������HY>���g�8|�ʤ�G0D�� ��z2���q!��PL�q&"O^(��J�+;�D�[2��,J�M��"O�y�f�k�^���N(X+���5"O����cL�u���F �L��"O���bM�IJ�\�$��(2����"O<���V0	W�X`'�  �X�"O]Ӵo��B|�D�B!!�Xxj�"O�`�#�!}"V��X5�-�R"O� 6�I�S��`@�­TzB`�"O@��6M��N�Ȝ(�"Jt� �"O쉒�AI:�0`ʑk̭
SΉ�3"O�l"���+,�,<���C�oDxtp�"O )���8R&*�hi)R5�"Od-Z�N`�H� 4)ȹ<6�\�G"O\ɣ7�<�<0Q��&���"O�0� �N9k���w��(k�b
"O��rC�9@
�5KB윣l��k�"O���F6)�@rd�	*�A�"Or0
rf� H��<��!	*5���7"O��  �U��<�P�m�:2Ż�"O8�Ԁӑ-�|풡�ћ&�b�AQ"O>���f�!�J�k�&��F���h�"O q��C�"�b�� ��#r��YY�"O^\jm�s|�� �P�$<j5á�'��'�V�ZD*�活%�ڵG�n ��'�l�!��Ӣ@�Hy��#E�2
�'�<9�#���Z��y!�"�2��	�'���V"�Hӷn�.N�P��'�(�o�*����d	�T����'�x�q'J�sy�@�#�� y��'� p�� �j2<��s���P8�	�'�4sC	x�NP�������'��:e��6M��� ��@dr�'(�\+�N�M0�:禚>'�f��	�'�:,!�!D�C� 4$]?�
aI<!��O�v�0(@3����P"���n�<)���D�܃�o!O���(i�<!��`�(�!_*����e�a�<)Q�Z�̲y�
��]Ԉ7n\y�<)�g,Nn<���ҭT<
��/�x�<�v��e�F�*��Af/�|3���<��Ƕ:�l0y6΁�{��C 2OȔ���IB~�h�!*��Dc�"O��a�I�o�� 6AH*3̲i��"O�
��B@�2L�WL19iZX�"O0l�e�&K.�<�@�J��qa�"O ��"�[*YQ>Xh��@�I�Ti�"O��ғ� S�hY�Ĉ���I3�"O����.2����E�t��ũ�"O�*%��Zf�!3坔o��P�&"O�T+n[�hAx1����LȂ8��"Ov��aGĒ8�hq���@ .��`�e"O"P ��O19s����N�.Mv���"O&Ef�ş�f�{�M]x�v5"O
�J�cKB��<2��F*<nd�+�"Obi�u��.�d:3�� �N��"OV�p�D�!�nd��IWH ����'���w� ��dޒ!����͸U�!��ZO�~L3D	/\����<�!򤑂Q��<;%�Y��hXdf�Nb!�P�N��'̀O @��/Y"9V!�$N#u�^�@���ޝY"�ȳ5f!��tN&�rgN�,Ί�0$�Q�f[!�dS�[�ba���p�h���"IZ!�� �3�钊� �``6ƽ�'"O<��@ۼ
k�paE͜r
0��"O�"��' [�5�Fn�b�Ĺ'"OJ�1��/_�`+��ɌM�@\(%"Oes%�-:+\d.K�T�:�7"O���ț�u��P�ȑZi�x"O���]�M��!#
$aR,�"O\!�DEL�(e�r�ԉy,�H�c"O0eYgc��Nb��F�.1��1�"O� ��
�(�ڴp�噠a-��0"O��E	ͫDT�WR2$4Y�"O����`[�SF$�Rj "Ip�"Ou���˧'P<��R$I��
`"O�Ufȇ@f�a�W�q�n"O�I2�BYW���8�$�P�"Oa�)�)mޮ�����=K�R� e"O��v�¹�H)��3E�0�:�"OȰc�NՋ:f�����J���i""O�Y��k�(0)��`�-�ЈP�"O�����I��!��@�����"O�Hh& 7]�x�ʜ?u�!*�"O6�3w��6.�ȓ��:;O<�"O*T����&�pq�rmM��y�"O��$U:' ~���֪�Ԉc�"O*-�e�^��AK�"z�J4��"O��C[S�������퐅"O��E�1Vh%8��Ne�^9�"O�@�/��t��y���7-?>�P%"O�i S�Y�#)z�c�$߷W!�]8B"O���r�H�mCiD:��A(�"O� ���,f�iQA�@����5"O���nW���:��N03�8��"OJ����( @S��/%��a"Oha $���!c��K!S	xU#�"OV!� �Fq4A��jPx�
�"O8���5i����`�[2p��L�"O
�RN�
<��=	�Z�r�.��@"O��UHD�-�P`�G\���B"O�U��o�a��Lr�`ȉ9˔i+4"O���W�)����`���Ñ"O���ChοKl��_�ay�%�"O
I��!0�1&��0w�X;�"O��)b��!"����;8���F"O�������h���� �X&ޡ�g"O>��Ǆ��<��dQ��lr�"OZ�Ři�
�P�ΐr��a{$"O��9��!zb��A�;r:P*�"O��	+�	�8)��@\5Al��H�"O0-z�� �D�Q�o��C0N��"O m��%�1�y�e�R0 (��"O����@�(��YS�AZ!� ��"OZ�91��o�� &�IP�q"O0ؐFO��&���Y�+F�diq"O�9��X\a��k�*A5��IB!"Oj!��.�t� 	�&
�s�^D��"O`�F8��#���"n�D"Oܝ�GA֙E=�8����C�jP �"O^�HvƐ��B�׳:�^P""O���P"�%X���A�z���xT"O6T���3��)���P��&�ȓ&����hǻz`=��K��>�>�����dJW�A�ϠD�-P�.'��ȓ]����6jװWt����H���8��ȓB�*��J�:?EKEc�����S�? �Y��\K�v��Ei��Q$h�"O��"D�!��M�f���+�D�P"O���q��8YB(�&�#=�j "O�a�c��80T^�qVV�su:��"O.�� ��t$Kwc�4VZ���"O��
WvB^��×C<�}bT"O��3� ٴ�Yp�S�u3�Y�"O��Ņ�0jF荙|%�܊B"O���I��n�5*C�%vz�`�"O�)8�(�*���j��]�"Op�`"�(4QĤzuL� �.�YV"O$�(�Z����3���r�d��5"O8q��l�F��=2�F�<��i1"OL�k�&M�p����&�1��m1@"O�����ɊhxDA���Ҹ�Җ"O�9�s��t�Y��Վ�x�kW"O�9 �N)8�y��V>�r��"O������K�$h ��.>޸)��"O$XhG�S�)�(��Řs�6E("Oj�q`g�$\�}�)�4C�a"O(Ȁ���;�p5C�fZ928��"O�] �A��J6�|J�$Ph* H�"O�=�Q��C���R�Y�yԝ+A"O���DG��^tB�I��d�!ұ"O���u��EܨA��G.xvQ��"O���q��0JG(�"��Ϗ*��@"O���3�M&���QX��"O����K�&��$��-S'2�6U3�"O8y��*X�`�ҍ_�RTp�"Od�fk2��@9Q.D�x�\@E"O~�:0
F�t�!A1�P�O�J�K�"OD��JϘJ�����6��MU"O�8[DA\�{���*�+�;-���r�"O���ň��w	�m�TK7u0���"OB�X��פHi�����]����"OƁY��ǿe���e�,W�H�"O��T/��&plx�%� �P� 6"O��������8Ѯ�w�nh�"O�"┆'L�*$D�$-��p"O�����=&��r��XP��("�"O���#tF9)%߂>>�ݚ�"O����H�4%���u)܍3$m��"O�,�S!�0N�A
���4�J���"O�".��S& (��^'xԆP��"OBXG��
=��#U�b���P�"O���wjQ=�L��B��l�~�Q"O&%&o��)�n����]�|���"O���gAR��iM;����"Or`��G-P�����b�T�n1yC"O����\,#�9��A8l���
3"O�쒠���M��+��-��m�a"Oژ�)=nhp����T�PH��"O�����7`���(f$an]	�"OLiaM;�P�(t�Z�w�4���"O�]sv�]�u���c��т��]:D"O|�u%J2l�T���W���j�"O���!	��_�T�pL��0x�"On�Y$� fp���9�lj4"OK�4�����,W�$�� ��y�(�73b������Q$F�jw�"�yro_��l����Y2F5�yc��:�yb.IS�|�z'hM�6�؍���V:�y2��&QE�I��^�.z�d�w\�y�3�82',�'1���w��y
� ��ǆ1b	� D��7�H��%"OP��<@��Db�i�J��Se"O2�bF��/)Ԫ����\bm"O�M9�lI,��a�"�	�JH:a"O��3j�-���cB�T��	�"O��:`�5k&y���9 m�"`"O���g��lpyKDkJ4
h�8"O���7
_9-�l-�5�7[Ӹ��r"O�X� �.=ԫ0eW"� ���"OZy��_���&��5�Ԁ��"O,��ϑ0Ő�7�2�A""O�Q�������٠�L��e!"O����MI7Z&���#ꃪ �(|��"O��25D/iS@éQ� ����V"O�)i��E7^�(-���h��;e"O��peb�թŉ�'`c��C"Ot� "�5}��`���}E��g"O!녉�P@R�ڤ��62��c"O���$�C�
:|X�'�sѤ	I&"O�e���]$8E���'�/��Y�w"O.�XS���5`�#�	;B<0[T"Op|�rG�^ך��o�W�Xw"O^ � H�5�*M�P'��p����"OZ�!+�m����ǵ��,�B"OF�!G�����wfτٖYr"OD��%g�F2���#E7z�P"O�Y��]�����5���˺�Y"Oz��%W6S(0x���:�L�X�"OD�[��܄0�"Ġ"�E�n�|`ht"O,葦k�.�Ʃ��`4-μ�h5"O��zQD�/N�j�� �S�^œ�"O����,/r�����f��F"O\�@�$%9��:�M�=�l0�"O�Y�C��,m�x�s��+:�>d`"O�Ī@ G"dB��Wⓣ'��A��"O:���'�usF��s"OFT���� G��!4E�uq�Y�a"O�q*e�<L�V��s����A{�"O�\K�K�1/ZR��Z�i�R�y4"O���N͑@.L��$����MH7"O��Y4↭,8B�aOR �b�{"Oje�R1���)�1Xrt	�"O¨��Sd"��{S�ɕpj��e"O�|�!.�̘��L�	,��F"O������I�"�UK�ibp"O����.F9G�5{#���-�ʐH""OL���b��e������5���B�"O�Iː
�	bdڷ�L��I �"O�� ���z\�BA�C����"O�!qO�H� 8X�j� ;��1"O�t�w��2q���cp�F�y���"O\}�gͅrl��(���;~�p��"O�p��-��#~���E��e���g"O6!� ��+@ t��%�)(u����"O =��/D1]��d$�*k�p��"Ovpu�VW�*���#PY��z�"O\�趢F�V�	�ĵL% ��"ORE�s)��:ϸ�#%�2K��z�"O����W�N,)�d�C��(sp"O�Y��_.Z@���;�l��"O�QY�AZ�^�����P�Tǂ5�2"Odx��a��2��L�6Űh�s"Od�j Ϲ��Yoމf�8�U"Oz���D�.i;R�	�h���	�"O� x�J��3e5�p
4�T�FjVus�"O���$"�
�p8�k�`\��0�"Of���J�޽(�䞛i@2g"O� ��A�7����iA�VZH�"O�͙ �K!��$�:6Gp��"O(�id�ؕkp�mH��k�B���"OT�I�W���H�#DN�l���"O���8N}\�2Fc���� P"OT�8�h�1n����@�À,"O:�pp��;�H��G�A;ь���"O&E*!���L�{� �p�8H�O\�
�,V�:�d="�lݜ  ��� �8D�T�22�28��qin�֭5D�P1�� q>��``�؅waFu�4D��k��S�Zk�H�+�h�"yꧏ3D���c�˛!n�;t�P�9O�\��C7D���OH�N��䙨k���06D�d� A(�BH��b�.,�袦�5�O$�	�Б�g�f���S��5B�6�=���D�OZ���W��XL���6�`�,D�����?� � ��	r�&T�6D�sR��:E,�ٳ'H�y�x���5D�ȩ�aL"Ἐ@Q�]Ȅ>D��BqD������D�e���qv(;D����J_:k��	�T�УB�����#D����4�LP�U�ͬT^˥f�O�C�	�$V��8��{��C'��"��C��,�N��'g�%W��H�ȟcf�B�I{H��g(ǎ>
!��+�-9]lB�Ƀh���z`뛍���Ha.j�`B��4j�u�̋f�iP�	&���[�p·K�CҶ1 3��Ԇ��
% Q��S�"�
K�p�y�'�a~Roɴ*{�M:c��0�$m�>�y��ė$�|!jR��T�D�&�
-�y���8�ҭ���9t0( 6lͦ�y"��6
#�<�V�L�Z�D˶%�3�yr'�gi�t�W��/O��Qd�?��'nz�2��B=$
�괤�F���'Mx��Õ�0��9٤��

,�4��'��]�0�O�;� P��G��}�V� 	�'Wnh�"�5A:��w��t@����'�.	�d��� WG;h'���'����!���A��IC����'�z@��퓄'"ݘA�+龠�.O��d-�Sܧ\	иZ��_isxL�ө͸�r�E�R��ɱ(�"sQD+51��B�I]S8�r�j��` ���l޼
s�C�	�:^��'/�'*�pڐ
H��C�	�D0=(�AD(0i� y�ȯ �zC�IC�T|�"(�6�h����bC�	������QȤ�p��*�*˓�?���S�k��;#����1y�/ϨY��?��I��R]@=;C֕?�(�&G߄HR!�D�(HX��j�/�%����/@!�$��~F��#�����i�*�	}�!�Q3o�eX �O8e&�
����Dp!�ḏ5h�����0!�*�'�Z!�+pm�ٙ�ᜠm��Z��գ;;�"4O�`��D	�� Z�_�[��8�"O~@��h[�=+��R�J�|��EX�"O�93q�(��5�4��x�Du#�"O�"胗V\m�k�Fђ"Oرd��>}���Sge�j�v��"O� R@��E�N����1��x�<!I�"O�I��C	�6�L��&�W�@!�@"O���D�;m��x0%��XѾX�Z���'�2]��G���՝J��C�����=JVO��'�ў�O��𱕊?T��Q��YX~}��'��L�a,��֡{�C!FF^��	�'c�|h�~TA���DH��'a>-RQぱ:��� �/A# ��
�'zy�U�*�"� 1N:���	�'\��V�х/�!"�d�>I�p� ��d�<щ��g��<��K�&���"G��C�'�ў�>�Ri�8d��7d��0�!2D���ԧZ�{zzlb���-�b��$D���d�X.0�\m��I�e�L	�!D�(i0��:=i{R.�Uw`@)�a D��� ��K����E*	<�b7�?ړ�0|��@T�YV<��CII��I�!�vx�p�'@*5Yu�Q�@R^}p�o�#䆼x�'m���A]"�b��S�ȵ!YH��'�xZE�M=�$=�W���b��]�ʓ3~�œv1�����)A�y�ȓ��aN�`���Cə�{�\��KA�� �L�"3�y�b��|8��I�<)��ބ&�N$˱���U[>�y�ቚ6�Q��1F,�rT@\8X�TB��3�΀)EE�W!��Sg��,H3NB�ɝw��5�W
�?��Ͳ@�(FNtB䉽�N�(.�P��՚�.N� V�C�I	�|�a��G�p��C)�'6HC�		)�#�gL��X�bm
yn���o���h���S)S������66�I���l˓�0?�Ҥ���Ƞ��o��B�����Y�'�?�����A�Q�"�I$: �-"�*��'�O�̡K�.W7��#W �>w 8��"O�Lq�o��r �z�O�,!�0�Y�"O�Q8%o��e3f�ۢ(٠;*"�'"O�x�	5 ����c�0?�����'��O�⟤�	�<Q!�ͽt�b�ڧ�)�����F�<QFD}�9hA��XW^Q[��Ix� �'��	�Y8��#Fڇ-r�\�'���^ B�
[$�!yEE�p�*qZ&�����B�	�y���s4�D�r*1��ꁽ�lB�'"�����(g�����ýWY�C�	>�t��A��|�`N��:��C�	�7��K�Ʊ���#U+�pUB�	�4��zHJ�B�h�$ "(C�ɟ�,�x��7ZC4�VJ�t<B�I??5R�x$�"�rW	�gz�B�	�gT���g�^����ˠ5<zB䉬@����"U����Պ	|�B�a1d��{�����dN�nƂB�	_f����C\��d�k�-�Ά��Q4 ��@+ЂI���%�ֲv��H�ȓ]��poM5U����B�91�H���}�u��jZEL���,E9-b̈́ȓ#�EM�_0,��Y�Q�E��x��pHƿM��#�Țq��$��et6���a[j��5+���nI�ȓ��4!�+�9tT�0;�暐Whi��O�,��/�
�N�G�P�kJ�-�ȓ+'�A*).V���t"�k��ȓz�-:g�D�:#Jx#'=FZa�ȓv�&��SB�=D\,X�c�ra��ȓtV� B'��n�t��%�0wҩ��S�? ��
��+6��:#�9��p��|��'U�-�mO3[�(3'�F�AB|P9+On�=�������xq,Һ�$X�P�F|+ў���I�.P�B�o�!]*��� D�$�PC�IPe�8:7�Ρ5�|�*�M�)�C�v�HՉ�e�-4�
�a�
x�C��&�P� �
��-�$�^�^��B�	�MҘB�
a���@TF4h ���0?I���v"(@h%��>X�P�e�T�<�C�1Py��1f9k�9;1�ΟE{ʟdc�(�1C�2%lR[¯�#��%A�F&D���Rϛ<Y3x��4���̤kUO%D��ҡZ?T�AB&GP�e��X��.D���2�Ծ0�H-�QΎ:=DN���%ړ�0<A���+�Z9@P�Œ7!�q�W�[qy�'m�`�ʍ{瘑x� ������'�XX(3e��\�p1�I3hd�����'��Ov���<�A쇫o��P�"�V� �(�sB�m�<	�f��6%D���b�] ��6*�m�<y������BL��
��BJ k�<i@��P�$b�B�^��8*�`�}�'�axCӠm��!���E=�@ek��y"oD��(5ra�ԙ>��qy$�D��hO���,�'
�����P';z�mY7G��+.�G{��'g�A4&ɛfJ� �3IZ�>Y���'�m�b�ǡn�h�#.2|���
�'�Ƭ��Oƽb�l���eЭ*�vh�'	�Ւ��kk�X2�(�.�{	�'�(�J��$|��|re�ڤwĠ�	�'Ʀ��l�Jud ��� i����>�'��	�µ�Ҋš���hU��ß�F{�����@�D��UK�����Ƥ���=D���1�H�*c�pѡ�1nh9e� D�Ի6o�_}�`8s�_�5\���H>D�4Tn^���Xk敒��:4��b�$�&�<�든�+(@��"Eu�<�bJ� 6H����ݤ3S�AXa)z�<���F|x���ȩfHnXJ�&VZ����<	���(]��"å=I�Ր��r�<)򁈼R��s�	SV.u���q�<�l�C#F@�)��fj��s�Q�<�D�4E���PU˂:J�$M�DO�<)��ʚu�E�v��Lp��6��H�<q!��1݌�q�n�*mUTQ�.�G�<�s��U�5�VdY$yﬀ�s��A�<qq�ð&Zdc��+�B���h�<qWk�l*���p�t���;/�Y�<6#��a'`�c�!ЄHB�4@��<)��܌w6�uRE
[=*BI��/y�<1Ɖ��"���A��p���	Dr�<YU��W�4�����˖$�s�<��lׯz���,�$<�t#m�<!E�N(S6 �mN `=�%�j�<���J�s���w�]a�^L9� �@�<	T͔"L_�D9V@F�`���ZG�<A!�O�)���2��A@%FuxO�E�<�7���SPFPgb�]\M��lT~�<�bGJՔ���9t���D�Rx�<Q7�Tl~D�����o�\M��/Rr�<��'I����h�Zh8���X�<u'O�}P3��@�n*Xq��U�<��=.�șz�T^�qqKx�<񃣒:FY�Q�4��.?���D>�D���b"C�R�,E ����d��S�? ����w$� ���nǺq��"O|�[RK���a#��N%|�j!9"O�8�4��wF52��.�-�"O�E*c�L�w�t��4o9F��"OT���O�H�\�s�n�i�RY`�"O�-)�̺I�
@aB��J-�U"O
���mT_�
���aڮD0�"O�驢���d�0�?Iɂ���"Opd s���?�&�����(u�'��	���(��U*!��E�T�N�F$�C��;Jd�Kd�E� v�ܙ��1Z<C䉭m�B�c��4'_� �����B�;[��!d�*i� ��"l݁d���0?���B3@��1�S(�?X꼱��_�<����6��i�d�ML�i!!c�W�<q�)���y��Ι:�~�kpJ��d̓2��(W%s���R�)�8ZR)��^(���K0��q"��Q-�T���=�Uk�]�6�
����g�u�ȓ"򀈷�) ��'��#P���%�؅�[�z(�f� K��ȣ���^j�C��9<���`%E9��@Ru��e��C䉅O��X��'^�Ĩ�7���r������/6�@ӕAF�7,|��w�Ɯ@w�C�G�V�p�⊽VGJ�s-F!L�B�I�f�r Q�T-�<5pS�+�\B�I�[-�1��߬+M$];�K�P2���O���D�. �r5�s!Y�T_�ܪ�?!��^I���h�I�2ET��I,��nq!��V���&Ý
~ ���L�cV�'R�O�"<)c��6f�`!���q��a��T�<A6��-Vh��@͉d*���b�g�<���p�N�ʐ \	;-�@4"Bd�<ɣ�<���.�j��Hu�<��m�=k/�	�a��0�J|���N\�<�o��!�LaB2�$�
���N�<�uL��&'�|�5�Q�rr��jC"�R��P�<i�K_T��ͳ��X�O��J���f�<���M*�D�E�"�8)���`�<�.Ҏ�McA�D8<��Ģ�A�'a��O�FK�1*���4ྕ6l�y��-x��'N:2�������yR��/VѶb�.U�;�\i"_�y�H^9	"�8�d͓1:��Л�y�B�7V�hu�䃏"8p�x7 ��y�$�5H���#m^����aMM��y¡�[;�E��Y�,"us �˓�hO��D5�{w�](����aHx���C�_4�]'�F{��DF΄z���6Y�
�����y"�W@���� �<�\!��?٘'p�H�M��P��
ߔ������hO?%�`	>2 �G�Q�%r� �8�$8�S�O�Hp��ĸ$�40�F��nx��"O�i7JŖELT�ek
�ba��r"O��Pw�K&!�i"�؋pF Y��"O��8�F,ZAc	Y(VA��"O$�y򎂓`ȀC�Ι	�L� �'��D%�, ����mx�rU��0z!�D�	<Ґ��V�
��"KHR�)��6)P��NA�>�0vkM��Q�'[:�S1!D�c�4��Ej!��Y�ߓɘ'XrMp���r\��Ĉ-�
0���?9���I@��*��v�S�t�>@�� --�C�}_ސk�#�5'�r���ـ[��C�)� ���AG$Xz�m��@^���24"O�ċ#隤*���k/]�_���;��:LO�����"<Yh���N�8��F"O�ViX'[�,hb��Gs" �P'�'�I
&h�仢�B�\��*���)O�B�IR`��q�@7!�>�⃺3��B�I#}݈��Q��Bi+p�F�+�B��+2��`��_12<z���PT���I^�'f?y���)�c�9&�*0j�)��0<�2'��a�X��UK��5t^)���VI�<�$o�n�xQ��N�?5�����Jx�t�'b$�	��M�<xhQ'*R�~���	�'m�$X4�A�U��8J�/��tn�T��'�l�GH�'hĐBBME�0�R�'��h�'E d4΅:Whӿ=�b��'���VD�!<l�����[���*�'bF���:�S��F�}�
�'-���U��s�`X R�S=-���Y�����*>�^�����5���:4e��!�d_2~�(�g�3x���y&*I+*�!��+Q�kK��G�F���d"Oh�pዄsl~�qufQ!�� �'���9Ll�y��L�iS����˲:LJC�I�ru��HW�Ϣ ���6��5�C�<p_��b6bߜd1��@�3���d�O�{�&�ZrkE-i��3��}Z���Da��*4l��7����J#>����7����
��e�*Q��6�XI��Ga(��RhX�	��Q(q�`�ȓh���9%n]+s�pu�cO�&4|��ȓ�~lA�AY�@e|�q��u���z�Լ	�� ~�7���t�ȓ4�䁈e�	���w��}N��ȓ\ddkBĔ�8����,DA�a��q,���.�T�! ���v��ȓB�|�ZG	:X8�(V�J hB��%��E{����
�N�8F)׈r����ڛ�y�N!����R��RJ�AX%&�!�y��ʅ �x���1=-�%C0����y�'��jmA�Aͮ2� y��c��y���-��	�gi�.*}��8�!�$ȝ4����#-Q,�Cَ�!� =NȆq!7�ЅV.��!!�P�!�d�
q;�;�7F�Ys�O4�!�#�2KL�w�Z{���ʠ"O�Pg�åe�d�"H��	0�����';�Y"?�`���V�@���!L��^y!�бp'b��"W!1N�j�+R8=�!����iEGIfpR0QQk$z�!���3c܀� ����mq5��	�!��|>6-�s'B�\t !$Jp�!�Q�k(�=�P��'{�9�D�$1�!�dJ�p��( `�B֚i��B�]y��d w{`*r�ʿ+�ށxv���~�ޒO����D-mܤ�׬��JSV;��E'NS!�+n�pƪA�S�0�:�cS%Yo!�H
m����SF�����ԠR[l!�Ӕg��*��ٸC�nM�Ϲo[!�dÙ>���H�j�ۓ�$;�E9�'Dhh�fN+B���R��=0xމ��'z�%k4�P�*�ȱ�E���$�F���'�x˴#�.}~��Cd����H�'�\ex���`>j9S��5d�0�'� �,��vA��j���^h���� <�Z��W�m�J�ې��QF\�W"O���A��QS������`�"O*|)%�/^8��_2�!�"O]�Ԭ�37���hp,�&|�I"O��@��6S��,�MB*&q���"O��� ���X����M�_Il)�"O�e�B�ʮB�q��#�98����'�'ў��J�'O�����-;�9�r�
�s���X	�'ZDѨ�oӳ0�N�j.A)��[	�'�~|P')�k��< ���6&����']<�U҆K��D��/��آ�'SJ�����g�`x��������'�I�F)1^�x-��J���*�'d-
��W�-�(2��IL����'�(���+M,^ S7��/q��	�'%(z��%/����v��8n9��'��}(�GĖ{�y��kщ����'yp�c�N1��	J�� *q�Z@i�'Y�\(Ӌׇb�p�b"C�}��� �'�;a�Q$yf��@��?r3���'۬��P`�;xe��	t�,g. Ě�'������Yb�y�é���z�B�'?ax�Aҭ\ x���6�~��K�"�y"��V����s)�dPvkB��yR�Nyr��w�[CZ�P6�� ��O��D�Ob>E`@����c��I;Iڼ\��-D���f�[��p �BՕʀdaB++D��)"�-2 :5���f�5��'D�h@e�ΔZ�>U"�ǥZ���!��O���!�O����-u[��yq�s4�<� "O���!m�N�f	��M��+��2�"OT��C��fi��	GoKZ	[r�'�"��|�K>����;x=mH���	s��d�2���'1ў�O�rȑ	T�)q�l9��җ'$V���'J�j	�al��C kݓp�6L��'�F��!	M��$��Ă�8�Rzyb�'��-rw�X*Ҍ�	D�[�>lƬ��'�T�uO(���X#��/%p�9��'t1��#<}�,h���2���/O�=����'B�a�̧y�(�a�ʣg��<����y���_���ёn�<0��%����y�� �m���/>F+�Y�y�IסCj`[#�U2IȢ�A0�y��Z&�j�8�FR*1n�$��n�yR*�40�}BӍ" ��:�� �y�H�/ն�ˍ:tZdjb�(�y��ޫ+&�Ȫ��N#�|S��y�`ٶf.V�33��.��$���d!�O����=n��A2��-4J���c�OE�@�2lؽE�R��͎#��� ���2O���cB�:�Ձ�n��^H��"O�ŊSfS�+_�݉ Ó	cb�L�d"O�����
+^%���
R��%�P�'�ў"~b��L�Q��}	)

 ւ�RC���yb̟0>%���/M�Ayã����0>	WF��Kh L�ä��&�(����c�<�V��^T�(�!t�@d��h�<ч˓�7��|�b�؅jK����N�<!��V�	H�����5U�l�A
J�<a�kN�t=��a�� Flq2id�h�?ɏ��Obu@�Ɖ��ۅL�7  �"O �2i۔:�yxD�J1c7�|�'(az⩕kz��&�J2[����]�y�nä!�L��C�;�M�cOϴE�!�� "U�F�2UV\�3A2g��q �"O؉Sbc�J�@��]7��t��"O(8�rk�x��J-ٜ~�"u�"O�����@Z؉ �f�"z��H"OJ2 g�*TJFf�f�J|{�"OZMz#�E9	T ⪈�7!�E�P"O�HS*OoP���IƦ6��"O�tK��;h��8�C�4`��V"On@��ƕpf:�b�?VQ��q"Oƀ9����]
��'��@��9��"O���E�b�B(��c�V�b髃"O^�b��J37�~u�s���B�TYS�"Odyڄ�׾?�,��
��h� "O&�{t;xXp��jЭU9����'��'�az����<8�P�$D@�6���$�G��Py�(��C2m�����W@M���m�<1Tn�'9۬@��C�\T,}Q�,�C�<���ǨvitL��� �|i#�Dz�<��(����.�
$�<m*T l�<� H�1R��%���%)R\C��$Љ�3�=`y¯ӫ��B�	��捂�h�H<�i��-M�nY�B�I8)�T���`UP��Z��9!򤝁2T41�#��"��`(��@��!�DF�X�nq��-I! ��˵#7aR!�o��y�DJƆ%���P ��8!�d�*b����K3b��L q�-%!�D��h�L�)5�F.�d�m�*!�*xz�"r�`F����bN�On!���4%�7�. ݘ��_�GF!�&̴QaD�y�AK��<F�!��J� ��V����\�r��zn!���h�jLb��A�$(��}S!�dK�q��o7�N��deW�PX�	w��(�� ����:�@	���
K����"O�]��j[;�<���Dp��Db"O�m)�h���9ò��i����"O�p{eG�)��%�@�P�B��y �"O����ű+��Mqe�H�-�ޥ��"O�`Q�ō]�ݘ/[�B��8��"O��s���6����L�`��"O�TH�.tu�\''�R�X"O��DEӘ:(��e�\]x�CP"O�!ې�ˋ?�U���9R_ԛp"O$��������� �;-H ��O�(q�&��U����%HA�U}H���0D�t7@�;��d+�h�Z,F��).D��Rl��-7��D��U�8���+D�H`��ؕ�  DcQ,k��4!�H)D��)���+S��BM�a�l"!5D���v�P� K��S+S�HQ��6D��g�N�B�q�Iҿx ��;GO44�d`�(G�a�BP	�B[�D�h��OI@�<1��L|���������g�~�<�E��HGąq�*s�La٣OR�<yag�8AbU�'�!x����r�Kz�<%�F��p�u�ޞ<�hL�BGw�<9��4��(��M�'����wiK�<��@Vn�,1�-͂sr�5��I�<qrhJ-S��*`$����%kED�J���O�&̠P*�)H$z�	3憶� D��'w��+�	;/��E�k�Dyh�'�-�p/SE�h Ϙg��Qy�'[2��⋪R�p�AQ��6�A ��� 
�[c�:j}i0��F~B���"O��R�/;C���g�@�__��!"O�`�C*� a�(l*$(�6C��P�"O���kܡ	��tR��*G��!"Op��5��F&��#�B��M��v"O\yy�j%Ybj5�jM
�� �W"O��1�.1�����G*?���0u"O�]���{�f@x�Շ7��rb"Onxrp�SuO�����[�),�B"O��¾h\豉�H�9BF ��E"O�1�e��"��`'Nx0"O�\�FŖ�-DR�qbE;OtS�"O�����ք0H��B���n�"O��� �5I��	��]lޖl�"O�i�$�%;�TPi���^y�鸴"O�����p@��0�����yb�;S�Ĥ�!U�E��e"#�8��O�#~�F��+ .�&��>Q\�#2E�I�<ɣk�6]�갂&a��_�|��G/�n�<ib�ΜS��]BQ�D D�j���^h�<�p��$���# �� ��nK�<�Rd�:&妠y������H�C�<�����t�)uBU�T�8�OF@�<�r�^!r!\�"�(�[`�Q�5����#��'�(y�8۲J��J'��ȓE�(�3cb� }���A%��	dB��wP�dN��}�@�a�lą���`��ł ��Li���&.��ͅȓ�����Z)}���w�;>%��ȓP:Z���%Q�?��9��4 �	��V�����L2p�P�#�.�/z܅�x�z}����+�h�y���Q&�ȓeX���MS
i7�A5"E�le���ȓK3�Y�J�g�zݘ�D�$4��-��C \�؜B����F��Y4�h��@��%�5�7	F����S\L���'
d��AQ���)�g��C��8��1ib���sG�ȉ
�C�I�	��a��"����� >ա�d@�B��)S��9ˑH�?A�!�Ǉe�UZ�Q�	rZ��Cj��!��.�^|�P���DI��P���!�䄩�¥�㔐;=B�Iܚ8�!�oE�1`���WT�T�$h] [��}"��`z��T춑�!��t-��8D��*�ʊ�?��PB���,��!b�:D�L�f֚ cz�
�kZ�4=h��I<D�|`�����8c����~XF�t�,D�Pp����B�J�����3.���L+D�d���P����@��]��ɓ��<D�Xɲ�Gb��I��E8v��5J;D�42�+M9!8�E؉RY�P�3D�`��d�����,2��H`�2D��ʐj�AyL�#0�CRwx����>D��� ��%{f�f��{�)#?D�Ljꏁs=�5(�P���t���(D�XI�C�M(]ra��8{��bV�*D��$����b�@G�d���'D��`%��
X	n4IE�&�n<Y�d$D����!C�{MT) '܉%n�b�"D�xȦ���V�ڭ��I� e@���b5D����J��lO,0�a���.�Jp#�� D������I��0��n^�"*D��#� �7Qr�D�&ExS&Q[��)D�� �}���43 �ӧK�:Fﺵ�P"O)0U�K���t��[I��L�g"Oށp2��;WP9�vɔ�pk��A�"O��RR%UU�T�1��5�8�kw"O��!W�S�/�n����� $�%a"Ot�
R �F#R�i�j9�k�"O~A:cF b'*��Щ��<�b�"O�ܳ��N��/Ɛ#��iE"Oz�RB�I��9bV &��ݚ�"O��	�Ul=)�/�>aG��z�"OVI��J�_P��#�ͣ6����"OH�OIAnV��EL�5����"OdԱt������g�U<:X�P�"O-HP�\.mp�M0��V�J��T@$"Ol�GF��G���b�ϳ.���ip"Oz)�Q��9�Љ'�?��4r'"O���p��I_�aR̀Z��Ұ"O�A��K��Y�hs��]@��Ũd"O
��6dզ_ɸ�Z��~��$	a"O�Ջ��U�eY��FW���k3"OXz�) �$!� /���3"O급��o1�i�qj�
N@t�'"OH��s�K�d����#� H�E 0"O�H�d��--��qwc͗'�v!�"Oڽ�"E��My%�#� �g�$D��XP+����P8Q+��>i�܊�.D���&��8.�M�t3�KҦ+D�XebKN�jU
R�ޒI�d���#D�$"b)�2=�d�&,����P���!D����z����V��0EJb����?D���ЪD�YxFD�5��:�@Հ0D�d;g�Ƣ��� I/`�	Ъ/D�l20)���a�t#�j�M!��9D�� g�T3C�tY@OI�N���1D��q��;B�p��d��f՘����.D�*��U�ԡqv��n�8(�1D�D��DިX"��DBF���� .D�@Ar"�-i)&�7m�t���zą'D�(K���0��p��*Fd���'+D���j��T�D`%d�#":<iD�*D���gx���G�K� @aנ#D� ��i�s�l�)��ّ$�Hi�. D�`����R�Ji���ʦF�Tດ ,D�\���}]�щeȍ��v�r�+D�@����5
�Y���l1�GB*D��X6f�+l�����& T�#D�p�HǙ�H8b%��4�>�pL!D�LJ҄�kj�8�	_�jE�?D��X�Cзk���r���aτ}�T@?D��	�g�*(%���<�z�P���yb+��N�jB�ݰZ��a��y�mעE�&�!d"i�PڤaC-�y"��(�d��ʏ
x�IQd��y"���,x1����/7�r����ybo�i����蘤ĎQZb��5�y�k�R�<c�F�}H�M�A��y�mV'(:\�pL
?�@���ȏ�y�n�!>���qBրiϰ����yb�M�:�@����]�<���yR�S%��0�`�"T�ԱI��ݼ�y���;� ���hO�NNtl���R��y�C�������@���w���y��C�Gn�PD�"cX"'&Y+�y�E�nJ<p)���rYБ��N�y
� V���F��q#�Q��NI�c�(s�"O���5�!b�X`T�\���Ys�"O��"���+U�*�)�b��5�"O��� �Y�4�n�3���,���K�"O^��)	�>!tt�d��"e��"Oْ���T0Ĩ���Ȕ$��q"O l@3�K?H����9w�4��F�s�<iD�#���!��C�B d*�OW�<RK YƒѫRlx���`��~�<�b�S�'b@����uz��c��P{�<!p��jdbyv#@h�H�&Xy�<Y��T�B��i�+P��E0$��r�<Q T�e�ry�Q�C���X��/d�<�lBF��}IT�b�����c�Y�<!��˷��q3��V�(S�KS�<y�B߅E�X���.޻7r��
VFj�<Q���A��P0�V+�m�.]]�<	0.B
D۰i��-K�lv��KU�<����c� �� EkG�]�!�T�<1�g�R4�K�I��ʭ3#�V�<���5#|��s��
u��~�<Ie`�=�>Ɂtg��=�L���C|�<ɤ����0�6��:�݁�z�<��
��e?��A���G.��A�@u�<�e�?/M���O�b"�D���y�<���ʪ�5!��06��uJ�w�<��+��x2�h���y�X��3hs�<AV���$y��b�ÁK���ɂJ�I�<!�"�{��Pw��&�EO@�<���U1L�Rа�$H�7�)W��S�<���%��|Ӱ��4G�h�q�L�e�<�*A�|��z��JHV��d�d�<�Ї_&����h#T���+�b�<�p�ݖ=(��1!.[����Ty�<a)ۂ �@T�V�@46\4�"䀛v�<єN�rGv�R�g����R���z�<u��cLf%7A̹4Q3#+x�<ɧ�ڐ1](�����k�R�"~�<q�CH�Q-[�iD� hU�y�<��"_7K����J�0^�ĳs`�q�<�q$^(C�P]��&,'��VJ�m�<!w	�;=(ҵ	s��q����F�k�<!��Y�䈒`�${��ä`�<)����G|x���#X���s��NU�<�� Zq����'�'9�| ˶
 N�<��,=�.����čF:�b��G�<�j�	(8��]�M�4�j��|�<6���,M�\��8d��)���v�<�E��q��Q�gU6B�t����Io�<��G�5��	��95$<��W�<A�׹�v�P�e�87�f�P��i�<�d��Fܬ���߷������}�<��@�0tn�첐�]4s���sB+�_�<A��ֽa�u#��I�^D$�;N�W�<G�l��)��ލN^�L[��[S�<�F�D�Ŕy#狐�"�Nq:�u�<�'�P�/H<Iu�M�P����q&I�<�d:)��-"��P>)��KJ�y�<�RG�>:+ ��f�Xą�g�x�<� ��O!���3B�<N� $�BAm�<A"�";R&�P�߾(�J��e_�<!G,+���K�ü��@�#��R�<1S�ˮQ�:d�ů$��()��)D��ZC�C~X�Y�С��ҡ3�&D�� %�Tb�!�eB�OZ%��P�"O&@�l�/����&8&�P�0"O�
�k��;�@�t�boma"O�SIW'@l���C�\(d9���"O��r'&���}�'K$K "��"O����3�0�!�ڬp
v�Pp"O�� u��L���j�W��y�"Of��/A3t����nʲ���"O�0ആP�1" �2W���p�`�"O��� @�,"�z�ȁ��'�� "O���Ǐ�7��D��+���[a"O��!�#7�+I
	�^%��IUP�<�6��~\��҉A�൛��PV�<9�j�)S,r������AʘS�<�&㚬w��\����6��P��BO�<����6L��@ຣ��^�_`.���C�Qs@E)b:�)��-8���%�&�s�D�g��Ļ���U B�I;-���8jZ�A��d��Y�9B�I� rx�B�E@
c��R�;��B��N�XL��9qj~�3����2��C�Im&mb���@@X��K�@��B�� ���� �6u�8	�*�g�C��2�)�N � ��� Fڧ^�C�&Z欑8B�_�sB�d)p��&��C�	�}��`����R������)�bC�	�<�b�{G`ҟqd`��2Đ0�8C�	�k�lk�"	�#�j���*C�*�C䉈~��a�t�E4�:=B�BxO�C�I�:�H�c��Eo ]�t�A�0�C�	�%���ru�_e�(��A�b0�C��3 ���΅��A��^p�'������J/G�*d�
>s����'D:�ʁ+q���Q�jd��	�'����/v�tq�ň�f����'�l�ۂ��`��Qڴ!TV#!��'�D*d��`�*��	�G@b��'u6H��@H#%L��`��A�.���'�:��T����F�P�k���'U�U���ŗnGXh�e\�`�:�'�n�ԃZy��(��%���&���'l¹ʗŏ+Sh(��kP�l�ԼQ�'�������5��x�g�7a�(��'!n�Qu	̾zj����K�\�	�'�����9<�(�b�l	1VJ^(8�'� ���бM�r ��L(Hy.I�'a������Z�����l�>F|�Y���d؋�������K�XE*3c�6`6�I�"O�T��kR���Rq� �"O�фKY?x����4,GԱ�1�'�qO�Ȳ0��}�b�r��ۺ^�v��c"O������"�=	�V�"O�yaDÓ����X�}j:&"O��
��E�]���7���K��'�VQ&��*ǫ����X���'>	���%D�X�'�U,Iöq� ,6�E�«'��f����7*�y��=(e�Q���Yh@��d�<	�O���D�	c�ʼ��iώD��}yd�'�ў"~�����tj�����C�x����k���y� �F�1HD�Dr�-s��Υ�yR ��F	�yãm
EKr� ���{�����I�1(����
���eX�d%v��%"O�Mq�)�23�\HU��A	���`�O��Iv8�T�⁏"�j0r,�1��@1�7�O��
�O� �Q�����y�R)�j����Bv"O��C��Ԓ	�ڑZG@J�Yg���@"O`���C��b��crf=�ɓfFPH<A�GL�,y�%�7�ޟ I�m4��̦5�tW��'��ϸ'�ܠ#qiX�^C���3�[�\T@9	��y�DI%�Q��6ݼ�!U�5�y2�=�!K�D	<:1�!�������>)'��<ɒl6�Ve2��̖#CT�R6	N�<a�����уU�Q'n��1
���hO?�	�_��r��<�������wB�"�Iad��d���bJ�6-���(O��%ړ����*фn�����W�ww�ȓT�4���}/���R���i����>W�r��L���(�B:b&�h��o��D����:U) 0�"�E��,l$����	�-L��0䋇�fZ�ze�/6mR��$`�������K��Y�K
؎v�>D�|s3�؊{�x����N/E(td21O�O��=1����4�d�@i_tX1��a��s)�{��dM�Z�(M���y�A�SaX�v�If��H�Eص ^7 ���S�Bz�\��@]�8E{��Уn�2Q"#�͢{y<[�̛+6�!�� �~ċ�L�7
��q��߹m�'*�|be�-5��<�=T^��8��9��?u2O���� j������Ȣ	�s"O���l���.Ы�f��;�"	���Ie�OuH��ҁS��?^9)���N-�S���5����@�-Pr�R��=��B��H�$�����[�4��c�݅��:��/ʓ:��>�i`�:��M�O���t�������Ұ?���H3!�� 3�@�?
"�Mړ�s̓ʈO�OMц͗ ���6%�.�I{��i�ў"}���cL\�9
�>2[re�s�R�$e�G}���*#�� �i�+&�P��cH��`��G{J~��G�/>HPҊ�9QT])�Ri�<i&�Ϩ��&���qG�5Yg�ͥ��d%?�N<����!�$u�a�V�z��U'F(3���i�OɲE��˾�: ���O����<�ߓe.Zd�����:��`�R�bt�%��Zs�)�Ot��2��'��c2Ț�Ln�?a���J�b�שG1qfܨ�A�f!�D�*JО]Ç�]Nκ��G�M�l���w�d+}��iA a��hʶ(�&�@�a��43!��=S���kV*R ׺@�A�U:��O�'��ϸ'E��TI0�-��Hɻ}����Ot��,]n����S�4�b}y��@��$-|O��A�rh��=K�N�#��ǳ���	Fy��|��\�b�~�e��6i��]󥍐,�y K�j�	�%H*b�D�������$�S�O�ؘ���h�Դ�fB�T����y��'R�d���@��i�T�0S�:�'�����)1�A�s�N�I��h@
��ēn�6�y�LV�|�y��R�k��͓�~"��0�'#I�h����*	goI�P��<��'x�O1�T�J�Ú�A�����\��aG�����	�+F^�@��pڜ��V(_�I&���D �I�Eq��[��L(���؅HJ�1��B䉢Fͼ��#d�G��W��%q����dt��nZ3bXe����2V#Z���� 2JnB�I�Sw�Ixc��[�>}��d�5
�8B�	�&���"��HJO�m�a�<[@B�I5O�$�SQ�%-~"�f�E�2�$B䉳h� �q.D-,�(A�rJ:d��B䉮QQt���� 	���+u#�&��B�)� ������]�f�C'ʪ\��IN����*[f�8FǇ7S� [$�*?`�*�O��d�	�NI��s�^+V>L�aO��$�]�B�G�g�P��VL!�{���P> ���6n �-�ZtZ ],��ta�)_W�O������Vo�ͰV�@<�}�}B�~��#�����mO�ej����I����'ў"|�C'5DS��(���-9	���b��i�il�la�����*9~j�c��ʠ�ћ�@=;!�	���H8�`.|�9A�NY�ur�Z~�i
Q���'��zV�t�8��Wi�<��S�'^�Yׅ>R�ژ����<s����d��hYQ?���gZ�,��X�\&����W<D�X#b$ӈr�FihF�D�0&8h#����#F�)ڧ �#p��fS$��+̪a$ZŅ�	hy"�i��2�!��c��-j�,����iX��cVI(m|�ȓؔ*��̡��<}��:�O�(c��E� �0I���ƹq`>X��'�ʓ!�"�[�)^�e��C�ۮXP�d�'��(�Iw�'��t�Te�?�$U;dJ�
h��r�'v�r]SwJ��ë]	cM8`	�'`�yh�!��
a�O�0eў`�� @�$�<r�^([g�[~���7� �Bj(��D�Cmۯ8Ѯȇ�}ƍ��Ҝx �ЇmR5M��݅ȓ#��y`�)�0o�����o;��'��~⢂���p��n�9��x������>�J��iwHɫ\<0��LK�m8��4� D�(
�I�%�acRĆ�o<��S">D�`@V�א<F�9�F��9����h<D�x��ޕn#�����! Լ�G�W������
�@f0�b������%�.b!��̷0�LȢb��.�0j���OL!�!%�L�Z�'�S��8���,�!�d���ehsʓ�Q�bt
S�C�F�!���0;��ІI�R������!�D�?&�t{�E�12�@�!��7v�!�$C�u�60`� �$+ 	ᎏ<�!�Y�WG��R�Ll%.d�EY�q�!�V��B�ۓH��*�+Q9[�!�dY�=�1�W N�G�xu{�
�}�!�$�+�T�7�ЋUG���/M�!�DÓB� �ȅ���{:@|�!
��!� (Ӿ%�!څ%�d�g!���!�ؒkFV(�TG\�+�|y8���<"�!�:S6�M����^ނ�����x�!�D˱F���q�
�(y՘M���!��F6��6hL����SȄ��!��B���L�6�� 2�{@!�$��S�*��P�Ö%�(	����
/!�ݼٞ�k�L\�s�ു�*EnK!򤑈f���jfD�1s&�{��0:R!�䀰�6���Қ��B/�]&!��L|Q���ɾЎ<{��	[�!��'j��4����ܰ�C�;�!�D1�\�h�b�2�vp�֥5�!�䔃V�����iJ�����F.4�!�W� ,Æ�	N��cC�C�F�!�$��}��I��(]��
(#!%�?!�䗫�N�9B(��jBL@��!��)l��{2�ߺz>"�hP@\j7!�69��Yi6+�3#)L�1#��6!�D�� ���U�
 �c����G!�D.na���S1�0s.��u7!�� ��`�]���`/�
Lڸ��t"O���㓕1�ꑪGN� Ϧ�D"O�-�j�0)��L��x�D��3"O�栔�R!��S���>ΐ��"O�5�C@F�d	
 r �
PV4@�"O*�k���(<PafG1Y;NQb2"O��[ώ/�ʌ0bEB?kƔ0p"O���Vo�"*�L��F��Q�^5�1"On�i�-�~��AIV3y�r	�@"O �{VM���C.�o�<A��"O����.�+ <���ң
GCP�"OX<��� ��H�2)����"O$���^I�6TxpV`��l:�"O������k:,��d+W�Y�w"O <�dܸIP� �C�S����5��<T�謉��0>Nر�� �U01Oj"��D�Y�������0�H��"O0���һ��i��!ɳ�"OR�#a��,SIP�v�Їp'�l" "O����G9����Eΰ> ��"O��{��[�$'�����#kY��x�"O.xQ�"D�C{����E�8K��J�"OP�x�Ħ�X�ț)�-��"OZ�0f�E2"�[��� �"O�E���R%�|YTd4����"O�s7�ɾ�̰J��P�$4>9�Q"O�5�Ra�T����I+ �!W"O�!('a����Hsb�G�Pl�#"O�雒I������h�ٺ"OQ�6�_#�B�I��/�6H��"O�t� ��]դ�� @�t�sR"O�0�k��/ݞi ��[�tˈ��"O�m�f���و��Wo�2B���8""O��(�I k�B}��.�(H�00u"OB��C��U:�[�0<n�"O�׏ X�T��,<l#j�*O��{�ɒ?�v�3��Z��i�	�'y���	A7>fPِ��P����'} (���_c�lz��E�8���i�'���eF�9�p@�ãڣ5PFi�
�'�0�#ɜ��5ȳ%:%�0L��'���"���o*���j�&�:\�'�Xܻ���a
��Oe�Vܨ�'�x�&�J>2M�Y��.sȨX�'L&�p�!_ ��$�'�����'�Ii��G�77�!�jD��05��'r~�ۃ���*	�"Q/&�N��'��U��.V%:-`� V&h��'��|���2{tbp�cF�h�Թ�'��xI�T��@P�c��\��5p�'��%��!i�nݰ�"�<R�
���'��'�ť
�,۵�б>��UR�'�vq7o�!H������H�-6�i�'K@�3ŉ�0��Y��G�>���	�'ߦ��T���� �" &O�$�*�"�'�6��NK�-n�}��l�0b��a�'�r����԰w���r薧iq���}�)�G�.�G�T��6T����
-V��V� ��y"�C)k���3��\.+��,���|W6��&�/�$��(��I5U��Ay�'�oV`�7햕3.�C��"Xa]��E�o`~9�`���.DY(֨ ��|�'՗K�u�S
�\���ȡ���0=9FET�s�x����� '`�B0��bM�;�e�5+7D�|	�9%R:ՙ6
E�EE�����1��5GB���3�9Q?�rպP�@�ib��_��F�!�� ����.oH�!�� $�<1b���7���J�pJ�j*�g~�I^����`�x2Q�֊Ŗ�yr�˴!��ف&��+5
�h!뛂We�PKb�m���I;R��p²�C��b�#�=$���̠S�~���g��~Ro�\�#4��F~>�p�G�'�yr%�@X~�a��T!4萀���'즑�P �P�E��T;:�b��p(Q,)�p�� ��;�y�
�fb�l�����z�����K��� F�Lf�d�	
>�Hh���⚩ h�ˇN�	��D��I�̓��''��r�ƐtELљԠ]=[\�aJ�r�4MK 0�=�c�E"�$�z��6Rb�D�]��$��-ԙE�U�'[8,��&��Dbv��%�X2�9�/O��A��:�`����"���2Ƈ�;4J�i�%a!��������B�~x�qT��2e����D�D&���&rD���ޣ"��,��(�����;D��S푞�J��XA�}R���'6�:�Q�w'����c�\�!�D�&1��ܐ�.[~F�)2B@i�旙>ĕ3kOH��s�,l�""�0on:5��&�/�@�$"O*4���=<W� �ce�e9��ٲ^��RDМ,�`4�1�'Bh5���U#6���D�	�w$��u$�`��Ή/e5Ȩ�#!%�brF��,���0�,4�����}��\d�L!QLQ�2�!ғh
\p�uH<^x��?��".!�� 񁈆4L�� R)>D���̈́�cɄ�� ��"t�<ْ`~Ӧ��Ҭ�JDA��N�&Y�G�ܴ5��eHe�
0�9v@�|m���!(�F��U��`�1��zk��j@bj�̝aeJ�kFq���Zi���$��p��Y CȊ$DN\X��[�t��O:p���ޮ��'�<l��n�/z�$�i򃍒���6��
��uʃJ$9�4�'A��>ɗ�'&.>y�4�12�Hc"��~�tdB��3�H�}���DE'����Gj�D A�w�� �G���ع)�pȲp�'�a� @�#A���Q1NZ�k�r���.�>-:�H_��M�6��[�7�@�D��#��	�=X��ZLȂ�!�!t��z���l\�r&��<)e ��P^0���/{	�!�7�.U
�e ŕ>Q&�3����?e�D�3�\�R,�Xg��� <v㞤��Q��5��	�.Ա�!]�R�=:ɞ����C��5�'�"��4ʸFj[�?7�0�R�
"d�Y�H�`I�U>a80�L2W�z䙡U�PX�e��n?vI{�#�r��b)D�\Q���:�4*�&��
�d7��}P����!QlTa�@o�rUdTIH���|��F���K�,P�H�(�#��M�;�z�R,N�A)��D�<�3d�#d��t��-��,�w��=F�1JN>�W�D���d�tp���rMЃ@�$�*��M`�qOv{���1qE�����	�w�T� �A� /�>��e��b� �`�U
a~��Εd+���!@�Yv����a�Ha�By�ɫ�H��	�[ ���ĩ/����O���B��#ky���)�=k@����K*+�~�����л�1�X��E�	=�b5��j�4�̐��"f����M99ߴ�а�� ƖE���9��
z�0,�@	 �0D�,�.
*�]�'�8���гnY&|�W8F�TXBa� 64�A�ȓ=A�\�菾\���5�B�=�6�'~���7���8�D�,v<ڃ7��1��P�'�e�~p�����!��B�ɌKi(�q���Vxt��� C%��(xT��+�=Q��_8L�0�̓F�ҟ��B�A2��E�EM
Y�dE,!�`�`3�ַ)�axB�Ҧ-h�;O�]1wb_�#H����EA�7��R�!8 ä$����?�7�.`��3r*,O(�S���X�xa�%�$J�-QX�����V�/�<)��'�����)[�h�a�R$�d>9�2��!ͨ���Q.P�,R���O��(3��-K)>ѱ��t�� #�ΟԚ��LAr�)�@�4V��x�$�.N.4ٱ�dp	B5�,-�Q�0�P�@��ȾO2e�S�'W&1����҅��0,���⩎����b��WM�][^)/�� �M�dM��x��]**��('��P�j��Bn�lia!��E�	s�'IN"�J�F�	#jIJ N	����+̮2�|�x3��p��� ��I
K���j�֏3���������Lo�~c���`b	)�4�q»p�z�'&� ��GD?��=��m�8��5���LsZ̓�n�]�����* H��q��ʞ�RU��h!P�l�0/PX�;

�,�z"Gסw<2�(�'�j�����Ewtj�cӍsJ�H2��d����n�'�4�]�r��q8S%��:��� T 
6+�$:��u#����8��'��eR@���E�c���)�%�؉���6� �QT#��0��1AB�]}�K�,��C:�yCi'�؍�'�'�
�y���2���B;O�>0d�����̒�xr� 6=�u����r�i����S�Xt����%jn�q��ɸ���Y�FT���G"�001���<	i��`Ȣ`$�G��'+B4��ӡXf���'۹,wbyr"Ţn����.h���'�")H,�f-S [n���V��8,utY*�w��	;2G^@�z���o¹��0��"v��`4)��=�(��	�`@>L�5e��$�\:���79,<�KT(C�[]6I3��wwz\�3B�=E�:t���5'�X�]�����4/�"	du�B���H�P��-˛[L�[���\X�4�f�Z0���!��is��U�5(�$����Z�rPY����:h"i��B�[K��ᇔ�lsԔ��&R6.�0���D�>��f��1��Y�F�U8h��!
��*&DC؍��
Qd��2D,6M�#t��A��AJ���(֣ɆQ�M�B5YM
�[�+9q��H�ȍ8z6d�5Dq�p�(�O�`�Ç�7\D�s�K'�I�_��1A��� $\8��@�z�ꍻ務Ӧ�2��
u��i��Y?v�dB�B�GE�DP�.�����C���*Y�T/|���C��9+$R��Jw���7M+?f
��,cP� g�4�]����r�E�s��Q8����DJ��YA�N-`V�����u��P�rwJ����?\�� �صV��LÏG�pf�:��'��\+�/G�qg�fU.��̸AF�F��<�q�I)ybvA���	�kp�Adi�2����V�R���1�F���X�&�V4eS�� ◝ ���X��+�ɝ!���H�0OhUc��I�(r�Zw8�$�)�^�0��`'KC�yB��W���"��
MU�T��E��{"��
YX%j ͈�1�C���򄁴!��,2s�ɖ�M�	E�/��֤Ch�=�҇���R3����i�C �|=�I�2�w�<�C�I�%���Ҍz��xP&.E��y"�Q-�"��GKLc�T���#Y^�D���ε8�w���j1+���Ha�=-i�I��'�l�	�I�>[�
�c�*�c����H�5������>v�6��	�y���	�~�?)Q�_�z�D�i��I�?`�����J؟�@"�Gm`�j`�N�0�^�f�]1byx����.P�*c��`8�X��,u�r�K�+7ޞ����+�ef�K�##j�R��ƬE=��df�*^(�0�ʨ+(�T`���y�!��K��P��ϞA�J��+���>zfQ���;:��p@���\'q(B!t�ԋ/Z�ɴoռ49!�d�8Y���0 B4r/�-y��!2-Ё���>Q�,[�Cg\�>�OD�p&��9}*ru B8�&]J�O&l�P`G1o�&�j�"ܖK�:@
�t��VK.L��MЄ(��!��8�d�ȓ7PV����֌m-@`��W���ȓԙX���"G�E��R�66��ȓIfh��ַh��<��k�7oexU��6��Q"m޲|��2b�,U�ܼ��l+LQt';h��1կ ɨ<��<�da���e�X8�@�������j�<�"gkT�� -r�U�~H��CФH3�E�x�8E ���|��q�ȓk �|hC^oN 4 G�ksfH��'�Hؓ*O���i�v� ���A�'�l[G%ūRj���4{@e��'�⼩V��n�h�pM
����
�'���Y�
Pi�-���Y�
!֠Y�'���c����H�K�F^�*�'���б�Q$5��ə�f�z���'M����/��]�@)׵r׶$x	�'�
D�C/�;
ZD�w˟n+l}��'EL芕���a��p�L;c�j��'q|�X�H�U2�D	U�#Q�8�K�'L^���!��oi�̚�B�0wb42�'|`����#�|�� ̤-|�d�
�'R�j6�Y�L%�W�������'���	�nEy��@�m��c�'Ό�JlG�"�yF�>pҔ=Q�'�N�3E�ښB ���_,]a�� �'�ث��_�;�H�d���T;PUZ�'"��+�cPLEl p4�xH(�a
�'	��ˑO�dÎu��%��'�xDѠ�Y[�ڴx��?XGR���'�Y)Չ� )7f!#��W��I��'Ҙ��1m�Q8����&E$5������� �в�f�r�\P���ް� 1:&"O*��r RC���k�*Ǆ;8 "O&5����S8��RC[00Z���"O@���\K��T�]���y��"O���X�p(p�BT4|TR���"OX��5c�L�V����'��1�"O�P�fE�y���zŀ�M�J੐"O�@4"�?i��b3�#�6��`"O�$��k܅)����$EU	T�Xm�G"OqҢ�A� ��=ᔯV��͠"OD��M�����*s�ȟg�b�"�"O���g�^}>Ias��j��""O���<FL�4#�kq�nA�7"O�p��/&�Hs�*]�1�f���"O���e��:U���)�{[x࠷"O���3�W)�y;!%���Lb�"Oҵ
E/�n��HYf�^�D�  �"O�i:�I�0F\`��B#յ=�F4a�"O�}�3^�/�n��tlJ&b4�91�"O�!��
mX|U�Č1m=��s�"OR�j��Cb\T�K7E?�X �"O�|�AJ�EL �k.L�e8�"O�T�Q��#-��ep�۠_t�""O~=�[h���LJ�O�X�{b�<e9!�d_�x&*iA����'8P��UKZ�|!���,H�$�T0\�"�h��H�!�$��*�}���)n���j���M�!��&�&hk4�[���x�2ƹ,�!�DUpܰ�Kb�u,��S�1	R!�ĕ$W7΁��t�\���V�|Z!�H�l�`�Ҭհ<�&�c�A6k!�ҢI������\)3�)��iE�	u!��H�2�X�At+�/���n�=v!�56� �k���IVN�	"&V�}|!��ڶ�`T��"H�t�E�.d!�d�$t�F��F��wiT�Yp
.Hm!�čO �łV�Rm�(�ZR�;Z!�,@��� �C)u�\�i��<_�!�ā�:��z��ܩ\6�qu�D�Lc!�\�J�bi�����q񗋙 o!��-R��|�0F�N	,�#��+�!���-���4��E�������?R�!�d�68@��0��U��+��(]�!�B8>���p���۠�q�膾�!�䐕\Nh
��*���E%�!�$æw��G���HgN@�w����!���'�J��w$�:fHq&*�_T!���$+?�xR��\�Z
�@��ȷ,�!���0�3�06֨x�膴F�!���&��]� ��Se��\<	�!򄄖
��i��SQ�g%ѕSf!�D�Z.��b�z�M!CdT]�!��>&ȴB�@� �J�#I!�K�%��S��+}��Cjw�!�à����CH��(H4�!���~�v�1E�#l�Z�����}�!� �4���aDP�G.�3d�)n)!�\w���%�+Vʥ�Ĥ��PyB�02����ԫF}~���C�	�y�8���V	\�~]��
AHE��T#�	�`.�'"�����I͞]"������sk"O�l���R�}1�tC�ӮW)�E6D��/(�$�@v�<�B��� �SFpR4#q��U�<	�&�F�s�I/��ʒ� ��y
ыĹu���� �3�k��=��)�!��D�q$�'�Ό��-�
Y$�0�O��3V�֒���0��*~l����\�00@F�U� ��rX&T��<aS��$yX� ��M#�'�u��E�� 2�0B͡?��q��)s�T���B{�*,(4�X�dXĽ��g�7Z(�'˺�+��D����94-�+���$I�s��6D��*RF�%씈��0uA�Df��/ b !9H9iS�|�M8y�8�Q�cҌZb�	��0=���]�f^	�į��K2FLU�Pp3m���nL�(7D��
���=�v���N�`�����2��0g���"��+2(Q?��`��6R^��ՠ� t�j0D�{T�X�d2صy�O���Aq��B��}j�>�v"Ba������Ҕ�P�� m&��u-�<s!��@�/��Y��ص��|�&	^x��2K���,����jqO����h!���KF��,g�@��Q�'�A�bk�;~�I�Ho
DK��M��G�:�v�<-@���0=a7�P%�� �%"�e��l��Bl�&٬}�0�=�I�-l����;�B(A'�1�܌��GC�{ǤY�Ɠj2��@Bېc/�	Yd�ɸ*�-Gz��4l~J��Hq�'(�9��	'�H�c�,q羅�ȓ5�XR@R>(t�Us#��+�v�n�I�x���O?hl�S��M�9`>�����+�}��PB�<�QCTc��@
���4q~�U�t�Wy}��!@0�����dx���p�ށ
�%㒊ٮuhƙr��:�OԘE���0`�;%%ݮfa,4r���w�^�;G�Д��x�N����j��_ZK�h�V��
�HORta��D�D!����#��*)Дz����ʞq��-�=�yR�ȽKX ��3��^��S�T��ٴz��h�1�',�6)!��
y5�?7M�z�؋�D��G�v�ȕ�['m\!�G�0��uڗ����];![�`�p *��Z�|P]�gJܷp�+.�����1�_�POR����*3�8!��<�I�"fZ�SU�d�!bP�{%��?Y<8+�Y�a���e�L�h�<�C29��	�'e�ts�h�'JIj�k�$g�����5�by&��	p�l���d��,d4d�ۄ�Ֆ5 �N�t@�'XEL�)���>\!�$B�#�֠d_�^P�}3����"�(��M�3D���5�6&U&�a���ʦ�yW�H?��b>-���]z�ae������r0\O\II�@ mm���'��IWkשKRH��&h���D� �q+7}R����@"�[��@2.�2��V���0���=� 'ך�V-*��?�'��I3Dj�k�@%�Ba\/@���o6E�N9��L4�OF	h�*�	!��a��P g>6�� .�q�F�82�>!u�|�ϋ,*���ɴ>�_E�8ɐ1��{;<Ћv�ƞIr!�	�5nxi�p� 5)L��E� O�xr�Ɩ�|y���r\z����g�d%���h�#"�E1؈q�D(�T��Q�>v4r��"�y��+Z��[)p�x`A+3]0����|RL����I3�XY��@�]���s�̜f��<C6�2X���xw��6.J��v�Dƴ�J��Z���l�$)a<��Ĕ�4�^�IF��H X��#�7�DM`3kU��7Ñ>�P
�Y��2H����q�޽y����v����9�l �Pf\���I�K�|�s��'k��R	زW9$�3�B8An��	�'
���!d�1t�].]#	�'t��FJ����`!*E� )�D���$�)l�2�Z+O�L����lJ�t��"'�,���0#�h!
�'y��R�B�.M�� �.�lk�Ova��Y�j���	2�^����g��w�D��G�%�4s�+�����s�X�#�$� q����Pf�<�E��:c���h��ҦHx=0�O�\*�Ŀ?YZ���i��P���%8&I,��s�M�W4���'-��%iBIo�,���U"���$�I�uf��r��i�Rs'H:M02��*.}N@a�foX�8{�j�4?fZ���N̯|P^1�T%�<a��޻2��YQ���O����M��P#���V	2}�%l�)zS^����ic���k�-E�*�e�%$�8.?k�@qC�YTY���������5�U9u�ھF>I�j�Yg�p!3a�T[���A�'��AV����EI�:@DI�E$�3Q��R��S�`B��!�1���L:�$SD�#!j	" ��>�Nd�dc��G�2V�?9��N�V�I%k @�&5`t���`�C���?1���&���!��O
�҉� �� �{ �i@f�v�%O,@�Y"#�f���F!h=�x���؟�[0�OBn�>qǁ�W&6q�#����Dx�*�Ly�EO�[w$lScA���a�.UN[�����OZ��B#��P�S@�[?`�~�3L �T8�HpBCE��}�G�.y�����'jI��ݮGR�<�)Bju)�&�U8��jdŊ�o�*���W��uG�Ut�M��m�$�(� �bmQEbG�ny�� �5eh��B1����<�ՠδgm��J�\&�II4�r�NQx�^��\I��(�䐠	�F/�����x�<0�N��u�@Ah�"ޜ�?���~ʒF�&���1,A=�ּ�E�@F�	�{p�A7K�X�$'�5�w�O�������
�FM�Ql�',�H��Ve[Z�T�{��T��.M��kԺ��As��~�C2	�Z���Iӻ~�,a�U)�v2�9��=O6�����^�"�9�㘳
�T���is>i���y��#ڈ����8��1��!�"�?1�mȩ/?Dp�#�]�ذ<q4��<fn�ꄜ`�`4���l�f��_(عz�'�M�Q8��@�MS��9R%�$�0����� p��ǧX�B�R�A���H�a!,OZ��#H֢
��4F��v��3&��",ߗ9`�:�"��)�%�G�ɀ*��U�Æ .q/�hʢKаx,��*O��������*$l2����Ns��#��x�4Y����7�I����g	uN�x���S�y��f�*�(���I	�i. �irɟ�>ܑ��KB�>����BBXyR�o��~�N/E�r/�GG���1ူ=�T�r��iB�yP5h	�3 4@6�])[��SuD��|�A��dq�p1��;�ƚ~bqa%'�#DP��Am��wf����<	7�חl�(S��.�T�G��B6zm�v!A
4�L���`$~���{Wo� s�e�9�3ɟ2q��Ѕ�i���"Gj��)�ܘp/H$g�v��	�)�Ԍ+ �Ȥ�?�q��,ty��j��HX0��9W�]T<J��P��,e�$�%�]pR�i�4,O�(���л\�$����ٙb�dAQ��Y�c�`IY�'l���Ý[y����YR\�b�
E�2DS�Ď$���$":ٰ5Y�' 8Qa��n�.dJ���V���>	H�4	��ۙ�?�d�ً2�#|���d�5(P�'HT�
��@K�<��-��&�W�È^�
=��n��^�)���L�g�M�Nx�R��0�@Uc�~B�	��Ra0�c�+R΢}�gC�/\�x�&b�=!�$�"��e�%n�f�&�3P���=&!�$��#	��Q7��A��ё#�]�$!�D� #��#�� k�� J��I��!�䋐A@�q(2���q�޸����!�Q@���ɒz �P4�.�!�ʚg�m�u�]NdYhAM�o�!�A&e��� � '@/�Tr�m� E�!�>L1��'K�x)�&+ g�!��b�ƹh�X<0ab���r�!�DT�J���@D��4u��$��նX!�ƈ1���ҫ�0!�rQe�]L!�D�2IS��#�Zrܵ���>:!�Ė�7m �Ȓ%�-6~X ��J!�dK�&���P�!�; D�4A���C�!򄑬Z* �����:5ƌ��-6^:!�6d�bxb`㚛�]a��ժ%!��;b�db��;f�����7R�!��S>z��H�m��n8���pq!�«{����w�M�ph�fdP�Yf!�d6Sg�=9��ȗ|3�!k�$�^s!�ּ?C��23�(-�B�w!���>(&�SE�M�cz0a��cQ!���/1V�ڇ��\m��4�ȡL!!���)N����؈_f��w�H�8!�$�;v� �@ޚ8Xl����X!��e��s�ϕ�B��E���^�@_!�U�C�j����O�v�<0���A"A�!�h$2����h��Z�&�+!���?)=+OK�z�jA�G��&!��aTp�{sʞ�g�:8B&o!��cx�\)�㖮�dY���*^P!�DM3��u�/)�f���Ϯ@e!�I�j�8�Ç�ЛA֔�j���B5!�$¨s�� B�L��C��L��ES�U!��މ4��qd֌I�,1�UC�!�Dv�)�UNJ-����L2!�Ą�ajnͳb�w���3��D4n�!�� <������tRB�Q�T3"OP�Kd��3�P`0#͒�i�T�k�"O
���ļ/���%ؐ|�ѰP"OPeS��-��<9�N1.�(�Ca"O��"0)�;=���2��(
o��;d"O���D��_V�	I���3+svy�"Ov ���ܣX���ꆉ�.�F�p�"O���'�m��M��ɠcF�s�"O:�����5�T�`�9e�Lң"O�遵���U%pI�@(��/GbMz�"O��+"K�"o	Fp �Z�=5d�{c"O	P��N(i�t@�@�W[n�F"Ox;Q`]�ڼXfТ.C��I�"O�a8#�ǝ~u,,+�$��S�� *�"O\1bD�׻9�}�gd� V�Qɐ"O�Kf�;߂��q��5pLHa@�"OF ��bǪ]Lt�y0BX+-���"O8YKS���3W�	�4bV��	B$"O���ę�xT����3>$��"O�0�d(�?��B"���3���f"ODL�2#L��Hh�\�FP*���"Oȕ��$۴:�d�R*����"OX�ʵ͚�G� b��Z=�rp+#�d��:�lLS�l�/[Բ��`ɡQ�1O>43��J�x��͓�-߫rي9RA"O��p��=>�5(���	�R��g"O&eas�ǜ#n@���F^�)��"OJ�ї�}�:=�V@�2lj:��V"Oj�A���{B*!zeL�-bH���"O��RK�B�m1$%�2Qde�3"O�����1*�v��dasd��K�"O𠺖��
��ʓ�^�I�1� "O�(p���$��iw��H��L �"O��R�o%KɖXZ�A�BO�=�y�@�3-g���G:@����r>�y�L�6_��bG3#ƶ��QɃ�y�똨B���i���R%L�;�+�4�y�/�`�]��N�TXd�am�.�y�?$�r�j�/ўL���o�+�y�	�S����ůD.���$KӇ�y"�ΆdY�B\78�jd�%��$�y�'��.]̓��(Y'�8zb��,Z��a���'u*���&�)�'.��q�@�f�D��Ó�b�6�#rI��"�A���~d�wA�3}J?͢���+m_LD�)oָ\�A��-��Qڤa��PL>���,h�H!�1K9�IQ�%?�� a�z̳J>E��� 1r�a*"j�x)Hp)2$ ��y��V�P$�qd3o\xȪ�!���y��Y3l����a���� �]#�yU��B8�v�Z"��+�P�yB�V�L @  �